magic
tech sky130A
magscale 1 2
timestamp 1755812063
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 14 280 119862 117552
<< metal2 >>
rect 32 115796 60 120000
rect 1320 119870 1348 120000
rect 1964 119870 1992 120000
rect 2608 119870 2636 120000
rect 3896 117156 3924 120000
rect 4540 117156 4568 120000
rect 5828 117156 5856 120000
rect 6472 116680 6500 120000
rect 7116 117292 7144 120000
rect 8404 117156 8432 120000
rect 9048 117292 9076 120000
rect 9692 116884 9720 120000
rect 10980 117428 11008 120000
rect 11624 117156 11652 120000
rect 12912 117156 12940 120000
rect 13556 116680 13584 120000
rect 14200 117156 14228 120000
rect 15488 116680 15516 120000
rect 16132 117292 16160 120000
rect 16776 117292 16804 120000
rect 18064 117156 18092 120000
rect 18708 117156 18736 120000
rect 19352 117292 19380 120000
rect 20640 117292 20668 120000
rect 21284 117156 21312 120000
rect 22572 116680 22600 120000
rect 23216 117292 23244 120000
rect 23860 116680 23888 120000
rect 25148 116884 25176 120000
rect 25792 117156 25820 120000
rect 26436 117156 26464 120000
rect 27724 117292 27752 120000
rect 28368 117156 28396 120000
rect 29656 116680 29684 120000
rect 30300 117428 30328 120000
rect 30944 117156 30972 120000
rect 32232 116884 32260 120000
rect 32876 117292 32904 120000
rect 33520 117156 33548 120000
rect 34808 117156 34836 120000
rect 35452 116680 35480 120000
rect 36096 117292 36124 120000
rect 37384 117156 37412 120000
rect 38028 117292 38056 120000
rect 39316 116680 39344 120000
rect 39960 117360 39988 120000
rect 40604 117156 40632 120000
rect 41892 117292 41920 120000
rect 42536 116884 42564 120000
rect 43180 117292 43208 120000
rect 44468 117292 44496 120000
rect 45112 117292 45140 120000
rect 46400 116884 46428 120000
rect 47044 117156 47072 120000
rect 47688 117156 47716 120000
rect 48976 117156 49004 120000
rect 49620 116680 49648 120000
rect 50264 118510 50292 120000
rect 51552 117292 51580 120000
rect 52196 116680 52224 120000
rect 52840 117292 52868 120000
rect 54128 117156 54156 120000
rect 54772 117292 54800 120000
rect 56060 116884 56088 120000
rect 56704 117156 56732 120000
rect 57348 117292 57376 120000
rect 58636 117292 58664 120000
rect 59280 117292 59308 120000
rect 59924 117292 59952 120000
rect 61212 117156 61240 120000
rect 61856 117292 61884 120000
rect 63144 117360 63172 120000
rect 63788 117156 63816 120000
rect 64432 116884 64460 120000
rect 65720 117292 65748 120000
rect 66364 117292 66392 120000
rect 67008 117292 67036 120000
rect 68296 117292 68324 120000
rect 68940 117292 68968 120000
rect 69584 117156 69612 120000
rect 70872 117156 70900 120000
rect 71516 117428 71544 120000
rect 72804 117156 72832 120000
rect 73448 116884 73476 120000
rect 74092 117292 74120 120000
rect 75380 117292 75408 120000
rect 76024 117156 76052 120000
rect 76668 117156 76696 120000
rect 77956 117156 77984 120000
rect 78600 117428 78628 120000
rect 79888 117156 79916 120000
rect 80532 117156 80560 120000
rect 81176 119870 81204 120000
rect 82464 117156 82492 120000
rect 83108 116680 83136 120000
rect 83752 117156 83780 120000
rect 85040 117292 85068 120000
rect 85684 117156 85712 120000
rect 86328 116680 86356 120000
rect 87616 117292 87644 120000
rect 88260 117428 88288 120000
rect 89548 117428 89576 120000
rect 90192 117292 90220 120000
rect 90836 117292 90864 120000
rect 92124 117292 92152 120000
rect 92768 117156 92796 120000
rect 93412 117156 93440 120000
rect 94700 117292 94728 120000
rect 95344 117156 95372 120000
rect 96632 117156 96660 120000
rect 97276 117156 97304 120000
rect 97920 117360 97948 120000
rect 99208 119870 99236 120000
rect 99852 117292 99880 120000
rect 100496 119870 100524 120000
rect 101784 117292 101812 120000
rect 102428 117156 102456 120000
rect 103072 116884 103100 120000
rect 104360 117292 104388 120000
rect 105004 117156 105032 120000
rect 106292 117292 106320 120000
rect 106936 117428 106964 120000
rect 107580 116884 107608 120000
rect 108868 117292 108896 120000
rect 109512 117156 109540 120000
rect 110156 117292 110184 120000
rect 111444 117156 111472 120000
rect 112088 117422 112116 120000
rect 113376 116680 113404 120000
rect 114020 117292 114048 120000
rect 114664 117156 114692 120000
rect 115952 117156 115980 120000
rect 116596 117292 116624 120000
rect 117240 117292 117268 120000
rect 118528 117428 118556 120000
rect 119172 115116 119200 120000
rect 119816 117360 119844 120000
rect 32 0 60 1232
rect 676 0 704 1300
rect 1320 0 1348 1170
rect 2608 0 2636 1170
rect 3252 0 3280 3000
rect 3896 0 3924 2252
rect 5184 0 5212 2252
rect 5828 0 5856 2796
rect 6472 0 6500 2252
rect 7760 0 7788 2320
rect 8404 0 8432 2252
rect 9692 0 9720 2252
rect 10336 0 10364 2388
rect 10980 0 11008 1170
rect 12268 0 12296 2388
rect 12912 0 12940 2796
rect 13556 0 13584 2320
rect 14844 0 14872 2388
rect 15488 0 15516 2252
rect 16776 0 16804 2388
rect 17420 0 17448 2320
rect 18064 0 18092 2388
rect 19352 0 19380 2796
rect 19996 0 20024 2252
rect 20640 0 20668 1170
rect 21928 0 21956 2320
rect 22572 0 22600 2388
rect 23216 0 23244 2796
rect 24504 0 24532 2252
rect 25148 0 25176 2252
rect 26436 0 26464 2796
rect 27080 0 27108 2252
rect 27724 0 27752 2252
rect 29012 0 29040 3000
rect 29656 0 29684 2320
rect 30300 0 30328 1170
rect 31588 0 31616 2252
rect 32232 0 32260 2252
rect 33520 0 33548 2388
rect 34164 0 34192 218
rect 34808 0 34836 2320
rect 36096 0 36124 2320
rect 36740 0 36768 2796
rect 37384 0 37412 2252
rect 38672 0 38700 2252
rect 39316 0 39344 2796
rect 39960 0 39988 2320
rect 41248 0 41276 2252
rect 41892 0 41920 2796
rect 43180 0 43208 2796
rect 43824 0 43852 2388
rect 44468 0 44496 2320
rect 45756 0 45784 2252
rect 46400 0 46428 2796
rect 47044 0 47072 2388
rect 48332 0 48360 2252
rect 48976 0 49004 2252
rect 50264 0 50292 1170
rect 50908 0 50936 3000
rect 51552 0 51580 2252
rect 52840 0 52868 2320
rect 53484 0 53512 218
rect 54128 0 54156 2388
rect 55416 0 55444 2258
rect 56060 0 56088 2796
rect 56704 0 56732 2252
rect 57992 0 58020 2388
rect 58636 0 58664 2252
rect 59924 0 59952 2796
rect 60568 0 60596 2320
rect 61212 0 61240 2388
rect 62500 0 62528 2252
rect 63144 0 63172 218
rect 63788 0 63816 2252
rect 65076 0 65104 2320
rect 65720 0 65748 218
rect 67008 0 67036 2252
rect 67652 0 67680 2252
rect 68296 0 68324 1300
rect 69584 0 69612 2388
rect 70228 0 70256 1170
rect 70872 0 70900 2252
rect 72160 0 72188 2252
rect 72804 0 72832 218
rect 73448 0 73476 2252
rect 74736 0 74764 2388
rect 75380 0 75408 2258
rect 76668 0 76696 2252
rect 77312 0 77340 2320
rect 77956 0 77984 348
rect 79244 0 79272 1164
rect 79888 0 79916 1170
rect 80532 0 80560 552
rect 81820 0 81848 490
rect 82464 0 82492 218
rect 83752 0 83780 2252
rect 84396 0 84424 2320
rect 85040 0 85068 688
rect 86328 0 86356 2796
rect 86972 0 87000 2320
rect 87616 0 87644 2388
rect 88904 0 88932 1300
rect 89548 0 89576 1170
rect 90192 0 90220 2796
rect 91480 0 91508 1300
rect 92124 0 92152 2796
rect 93412 0 93440 3000
rect 94056 0 94084 2252
rect 94700 0 94728 1300
rect 95988 0 96016 2252
rect 96632 0 96660 2252
rect 97276 0 97304 2252
rect 98564 0 98592 960
rect 99208 0 99236 1170
rect 100496 0 100524 218
rect 101140 0 101168 3000
rect 101784 0 101812 2320
rect 103072 0 103100 2252
rect 103716 0 103744 2252
rect 104360 0 104388 2320
rect 105648 0 105676 280
rect 106292 0 106320 2524
rect 106936 0 106964 3000
rect 108224 0 108252 1164
rect 108868 0 108896 218
rect 110156 0 110184 2320
rect 110800 0 110828 3000
rect 111444 0 111472 2320
rect 112732 0 112760 2388
rect 113376 0 113404 2320
rect 114020 0 114048 1300
rect 115308 0 115336 1028
rect 115952 0 115980 2524
rect 117240 0 117268 3408
rect 117884 0 117912 2796
rect 118528 0 118556 3884
rect 119816 0 119844 1300
<< obsm2 >>
rect 116 119814 1264 119965
rect 1404 119814 1908 119965
rect 2048 119814 2552 119965
rect 2692 119814 3840 119965
rect 116 117100 3840 119814
rect 3980 117100 4484 119965
rect 4624 117100 5772 119965
rect 5912 117100 6416 119965
rect 116 116624 6416 117100
rect 6556 117236 7060 119965
rect 7200 117236 8348 119965
rect 6556 117100 8348 117236
rect 8488 117236 8992 119965
rect 9132 117236 9636 119965
rect 8488 117100 9636 117236
rect 6556 116828 9636 117100
rect 9776 117372 10924 119965
rect 11064 117372 11568 119965
rect 9776 117100 11568 117372
rect 11708 117100 12856 119965
rect 12996 117100 13500 119965
rect 9776 116828 13500 117100
rect 6556 116624 13500 116828
rect 13640 117100 14144 119965
rect 14284 117100 15432 119965
rect 13640 116624 15432 117100
rect 15572 117236 16076 119965
rect 16216 117236 16720 119965
rect 16860 117236 18008 119965
rect 15572 117100 18008 117236
rect 18148 117100 18652 119965
rect 18792 117236 19296 119965
rect 19436 117236 20584 119965
rect 20724 117236 21228 119965
rect 18792 117100 21228 117236
rect 21368 117100 22516 119965
rect 15572 116624 22516 117100
rect 22656 117236 23160 119965
rect 23300 117236 23804 119965
rect 22656 116624 23804 117236
rect 23944 116828 25092 119965
rect 25232 117100 25736 119965
rect 25876 117100 26380 119965
rect 26520 117236 27668 119965
rect 27808 117236 28312 119965
rect 26520 117100 28312 117236
rect 28452 117100 29600 119965
rect 25232 116828 29600 117100
rect 23944 116624 29600 116828
rect 29740 117372 30244 119965
rect 30384 117372 30888 119965
rect 29740 117100 30888 117372
rect 31028 117100 32176 119965
rect 29740 116828 32176 117100
rect 32316 117236 32820 119965
rect 32960 117236 33464 119965
rect 32316 117100 33464 117236
rect 33604 117100 34752 119965
rect 34892 117100 35396 119965
rect 32316 116828 35396 117100
rect 29740 116624 35396 116828
rect 35536 117236 36040 119965
rect 36180 117236 37328 119965
rect 35536 117100 37328 117236
rect 37468 117236 37972 119965
rect 38112 117236 39260 119965
rect 37468 117100 39260 117236
rect 35536 116624 39260 117100
rect 39400 117304 39904 119965
rect 40044 117304 40548 119965
rect 39400 117100 40548 117304
rect 40688 117236 41836 119965
rect 41976 117236 42480 119965
rect 40688 117100 42480 117236
rect 39400 116828 42480 117100
rect 42620 117236 43124 119965
rect 43264 117236 44412 119965
rect 44552 117236 45056 119965
rect 45196 117236 46344 119965
rect 42620 116828 46344 117236
rect 46484 117100 46988 119965
rect 47128 117100 47632 119965
rect 47772 117100 48920 119965
rect 49060 117100 49564 119965
rect 46484 116828 49564 117100
rect 39400 116624 49564 116828
rect 49704 118454 50208 119965
rect 50348 118454 51496 119965
rect 49704 117236 51496 118454
rect 51636 117236 52140 119965
rect 49704 116624 52140 117236
rect 52280 117236 52784 119965
rect 52924 117236 54072 119965
rect 52280 117100 54072 117236
rect 54212 117236 54716 119965
rect 54856 117236 56004 119965
rect 54212 117100 56004 117236
rect 52280 116828 56004 117100
rect 56144 117100 56648 119965
rect 56788 117236 57292 119965
rect 57432 117236 58580 119965
rect 58720 117236 59224 119965
rect 59364 117236 59868 119965
rect 60008 117236 61156 119965
rect 56788 117100 61156 117236
rect 61296 117236 61800 119965
rect 61940 117304 63088 119965
rect 63228 117304 63732 119965
rect 61940 117236 63732 117304
rect 61296 117100 63732 117236
rect 63872 117100 64376 119965
rect 56144 116828 64376 117100
rect 64516 117236 65664 119965
rect 65804 117236 66308 119965
rect 66448 117236 66952 119965
rect 67092 117236 68240 119965
rect 68380 117236 68884 119965
rect 69024 117236 69528 119965
rect 64516 117100 69528 117236
rect 69668 117100 70816 119965
rect 70956 117372 71460 119965
rect 71600 117372 72748 119965
rect 70956 117100 72748 117372
rect 72888 117100 73392 119965
rect 64516 116828 73392 117100
rect 73532 117236 74036 119965
rect 74176 117236 75324 119965
rect 75464 117236 75968 119965
rect 73532 117100 75968 117236
rect 76108 117100 76612 119965
rect 76752 117100 77900 119965
rect 78040 117372 78544 119965
rect 78684 117372 79832 119965
rect 78040 117100 79832 117372
rect 79972 117100 80476 119965
rect 80616 119814 81120 119965
rect 81260 119814 82408 119965
rect 80616 117100 82408 119814
rect 82548 117100 83052 119965
rect 73532 116828 83052 117100
rect 52280 116624 83052 116828
rect 83192 117100 83696 119965
rect 83836 117236 84984 119965
rect 85124 117236 85628 119965
rect 83836 117100 85628 117236
rect 85768 117100 86272 119965
rect 83192 116624 86272 117100
rect 86412 117236 87560 119965
rect 87700 117372 88204 119965
rect 88344 117372 89492 119965
rect 89632 117372 90136 119965
rect 87700 117236 90136 117372
rect 90276 117236 90780 119965
rect 90920 117236 92068 119965
rect 92208 117236 92712 119965
rect 86412 117100 92712 117236
rect 92852 117100 93356 119965
rect 93496 117236 94644 119965
rect 94784 117236 95288 119965
rect 93496 117100 95288 117236
rect 95428 117100 96576 119965
rect 96716 117100 97220 119965
rect 97360 117304 97864 119965
rect 98004 119814 99152 119965
rect 99292 119814 99796 119965
rect 98004 117304 99796 119814
rect 97360 117236 99796 117304
rect 99936 119814 100440 119965
rect 100580 119814 101728 119965
rect 99936 117236 101728 119814
rect 101868 117236 102372 119965
rect 97360 117100 102372 117236
rect 102512 117100 103016 119965
rect 86412 116828 103016 117100
rect 103156 117236 104304 119965
rect 104444 117236 104948 119965
rect 103156 117100 104948 117236
rect 105088 117236 106236 119965
rect 106376 117372 106880 119965
rect 107020 117372 107524 119965
rect 106376 117236 107524 117372
rect 105088 117100 107524 117236
rect 103156 116828 107524 117100
rect 107664 117236 108812 119965
rect 108952 117236 109456 119965
rect 107664 117100 109456 117236
rect 109596 117236 110100 119965
rect 110240 117236 111388 119965
rect 109596 117100 111388 117236
rect 111528 117366 112032 119965
rect 112172 117366 113320 119965
rect 111528 117100 113320 117366
rect 107664 116828 113320 117100
rect 86412 116624 113320 116828
rect 113460 117236 113964 119965
rect 114104 117236 114608 119965
rect 113460 117100 114608 117236
rect 114748 117100 115896 119965
rect 116036 117236 116540 119965
rect 116680 117236 117184 119965
rect 117324 117372 118472 119965
rect 118612 117372 119116 119965
rect 117324 117236 119116 117372
rect 116036 117100 119116 117236
rect 113460 116624 119116 117100
rect 116 115740 119116 116624
rect 20 115060 119116 115740
rect 119256 117304 119760 119965
rect 119256 115060 119856 117304
rect 20 3940 119856 115060
rect 20 3464 118472 3940
rect 20 3056 117184 3464
rect 20 1356 3196 3056
rect 20 1288 620 1356
rect 116 31 620 1288
rect 760 1226 3196 1356
rect 760 31 1264 1226
rect 1404 31 2552 1226
rect 2692 31 3196 1226
rect 3336 2852 28956 3056
rect 3336 2308 5772 2852
rect 3336 31 3840 2308
rect 3980 31 5128 2308
rect 5268 31 5772 2308
rect 5912 2444 12856 2852
rect 5912 2376 10280 2444
rect 5912 2308 7704 2376
rect 5912 31 6416 2308
rect 6556 31 7704 2308
rect 7844 2308 10280 2376
rect 7844 31 8348 2308
rect 8488 31 9636 2308
rect 9776 31 10280 2308
rect 10420 1226 12212 2444
rect 10420 31 10924 1226
rect 11064 31 12212 1226
rect 12352 31 12856 2444
rect 12996 2444 19296 2852
rect 12996 2376 14788 2444
rect 12996 31 13500 2376
rect 13640 31 14788 2376
rect 14928 2308 16720 2444
rect 14928 31 15432 2308
rect 15572 31 16720 2308
rect 16860 2376 18008 2444
rect 16860 31 17364 2376
rect 17504 31 18008 2376
rect 18148 31 19296 2444
rect 19436 2444 23160 2852
rect 19436 2376 22516 2444
rect 19436 2308 21872 2376
rect 19436 31 19940 2308
rect 20080 1226 21872 2308
rect 20080 31 20584 1226
rect 20724 31 21872 1226
rect 22012 31 22516 2376
rect 22656 31 23160 2444
rect 23300 2308 26380 2852
rect 23300 31 24448 2308
rect 24588 31 25092 2308
rect 25232 31 26380 2308
rect 26520 2308 28956 2852
rect 26520 31 27024 2308
rect 27164 31 27668 2308
rect 27808 31 28956 2308
rect 29096 2852 50852 3056
rect 29096 2444 36684 2852
rect 29096 2376 33464 2444
rect 29096 31 29600 2376
rect 29740 2308 33464 2376
rect 29740 1226 31532 2308
rect 29740 31 30244 1226
rect 30384 31 31532 1226
rect 31672 31 32176 2308
rect 32316 31 33464 2308
rect 33604 2376 36684 2444
rect 33604 274 34752 2376
rect 33604 31 34108 274
rect 34248 31 34752 274
rect 34892 31 36040 2376
rect 36180 31 36684 2376
rect 36824 2308 39260 2852
rect 36824 31 37328 2308
rect 37468 31 38616 2308
rect 38756 31 39260 2308
rect 39400 2376 41836 2852
rect 39400 31 39904 2376
rect 40044 2308 41836 2376
rect 40044 31 41192 2308
rect 41332 31 41836 2308
rect 41976 31 43124 2852
rect 43264 2444 46344 2852
rect 43264 31 43768 2444
rect 43908 2376 46344 2444
rect 43908 31 44412 2376
rect 44552 2308 46344 2376
rect 44552 31 45700 2308
rect 45840 31 46344 2308
rect 46484 2444 50852 2852
rect 46484 31 46988 2444
rect 47128 2308 50852 2444
rect 47128 31 48276 2308
rect 48416 31 48920 2308
rect 49060 1226 50852 2308
rect 49060 31 50208 1226
rect 50348 31 50852 1226
rect 50992 2852 93356 3056
rect 50992 2444 56004 2852
rect 50992 2376 54072 2444
rect 50992 2308 52784 2376
rect 50992 31 51496 2308
rect 51636 31 52784 2308
rect 52924 274 54072 2376
rect 52924 31 53428 274
rect 53568 31 54072 274
rect 54212 2314 56004 2444
rect 54212 31 55360 2314
rect 55500 31 56004 2314
rect 56144 2444 59868 2852
rect 56144 2308 57936 2444
rect 56144 31 56648 2308
rect 56788 31 57936 2308
rect 58076 2308 59868 2444
rect 58076 31 58580 2308
rect 58720 31 59868 2308
rect 60008 2444 86272 2852
rect 60008 2376 61156 2444
rect 60008 31 60512 2376
rect 60652 31 61156 2376
rect 61296 2376 69528 2444
rect 61296 2308 65020 2376
rect 61296 31 62444 2308
rect 62584 274 63732 2308
rect 62584 31 63088 274
rect 63228 31 63732 274
rect 63872 31 65020 2308
rect 65160 2308 69528 2376
rect 65160 274 66952 2308
rect 65160 31 65664 274
rect 65804 31 66952 274
rect 67092 31 67596 2308
rect 67736 1356 69528 2308
rect 67736 31 68240 1356
rect 68380 31 69528 1356
rect 69668 2308 74680 2444
rect 69668 1226 70816 2308
rect 69668 31 70172 1226
rect 70312 31 70816 1226
rect 70956 31 72104 2308
rect 72244 274 73392 2308
rect 72244 31 72748 274
rect 72888 31 73392 274
rect 73532 31 74680 2308
rect 74820 2376 86272 2444
rect 74820 2314 77256 2376
rect 74820 31 75324 2314
rect 75464 2308 77256 2314
rect 75464 31 76612 2308
rect 76752 31 77256 2308
rect 77396 2308 84340 2376
rect 77396 1226 83696 2308
rect 77396 1220 79832 1226
rect 77396 404 79188 1220
rect 77396 31 77900 404
rect 78040 31 79188 404
rect 79328 31 79832 1220
rect 79972 608 83696 1226
rect 79972 31 80476 608
rect 80616 546 83696 608
rect 80616 31 81764 546
rect 81904 274 83696 546
rect 81904 31 82408 274
rect 82548 31 83696 274
rect 83836 31 84340 2308
rect 84480 744 86272 2376
rect 84480 31 84984 744
rect 85124 31 86272 744
rect 86412 2444 90136 2852
rect 86412 2376 87560 2444
rect 86412 31 86916 2376
rect 87056 31 87560 2376
rect 87700 1356 90136 2444
rect 87700 31 88848 1356
rect 88988 1226 90136 1356
rect 88988 31 89492 1226
rect 89632 31 90136 1226
rect 90276 1356 92068 2852
rect 90276 31 91424 1356
rect 91564 31 92068 1356
rect 92208 31 93356 2852
rect 93496 2308 101084 3056
rect 93496 31 94000 2308
rect 94140 1356 95932 2308
rect 94140 31 94644 1356
rect 94784 31 95932 1356
rect 96072 31 96576 2308
rect 96716 31 97220 2308
rect 97360 1226 101084 2308
rect 97360 1016 99152 1226
rect 97360 31 98508 1016
rect 98648 31 99152 1016
rect 99292 274 101084 1226
rect 99292 31 100440 274
rect 100580 31 101084 274
rect 101224 2580 106880 3056
rect 101224 2376 106236 2580
rect 101224 31 101728 2376
rect 101868 2308 104304 2376
rect 101868 31 103016 2308
rect 103156 31 103660 2308
rect 103800 31 104304 2308
rect 104444 336 106236 2376
rect 104444 31 105592 336
rect 105732 31 106236 336
rect 106376 31 106880 2580
rect 107020 2376 110744 3056
rect 107020 1220 110100 2376
rect 107020 31 108168 1220
rect 108308 274 110100 1220
rect 108308 31 108812 274
rect 108952 31 110100 274
rect 110240 31 110744 2376
rect 110884 2580 117184 3056
rect 110884 2444 115896 2580
rect 110884 2376 112676 2444
rect 110884 31 111388 2376
rect 111528 31 112676 2376
rect 112816 2376 115896 2444
rect 112816 31 113320 2376
rect 113460 1356 115896 2376
rect 113460 31 113964 1356
rect 114104 1084 115896 1356
rect 114104 31 115252 1084
rect 115392 31 115896 1084
rect 116036 31 117184 2580
rect 117324 2852 118472 3464
rect 117324 31 117828 2852
rect 117968 31 118472 2852
rect 118612 1356 119856 3940
rect 118612 31 119760 1356
<< metal3 >>
rect 0 119718 1398 119778
rect 0 119038 1490 119098
rect 117926 119038 120000 119098
rect 116270 118358 120000 118418
rect 0 117678 2226 117738
rect 0 116998 2778 117058
rect 117374 116998 120000 117058
rect 0 116318 846 116378
rect 117834 116318 120000 116378
rect 118110 115638 120000 115698
rect 0 114958 1858 115018
rect 0 114278 1306 114338
rect 117834 114278 120000 114338
rect 118110 113598 120000 113658
rect 0 112918 570 112978
rect 117834 112918 120000 112978
rect 0 112238 1306 112298
rect 0 111558 386 111618
rect 118110 111558 120000 111618
rect 117332 110878 120000 110938
rect 0 110198 754 110258
rect 0 109518 1306 109578
rect 118110 109518 120000 109578
rect 0 108838 1398 108898
rect 117926 108838 120000 108898
rect 118110 108158 120000 108218
rect 0 107478 1306 107538
rect 0 106798 846 106858
rect 117834 106798 120000 106858
rect 118110 106118 120000 106178
rect 0 105438 1490 105498
rect 117742 105438 120000 105498
rect 0 104758 754 104818
rect 0 104078 386 104138
rect 118110 104078 120000 104138
rect 117834 103398 120000 103458
rect 0 102718 1490 102778
rect 118110 102718 120000 102778
rect 0 102038 662 102098
rect 0 101358 1306 101418
rect 117834 101358 120000 101418
rect 118110 100678 120000 100738
rect 0 99998 1398 100058
rect 0 99318 1582 99378
rect 118110 99318 120000 99378
rect 0 98638 386 98698
rect 118202 98638 120000 98698
rect 117834 97958 120000 98018
rect 0 97278 386 97338
rect 0 96598 1490 96658
rect 117834 96598 120000 96658
rect 118110 95918 120000 95978
rect 0 95238 1122 95298
rect 117834 95238 120000 95298
rect 0 94558 386 94618
rect 0 93878 662 93938
rect 117098 93878 120000 93938
rect 116270 93198 120000 93258
rect 0 92518 386 92578
rect 0 91838 846 91898
rect 116914 91838 120000 91898
rect 0 91158 1398 91218
rect 118110 91158 120000 91218
rect 117834 90478 120000 90538
rect 0 89798 1490 89858
rect 0 89118 846 89178
rect 117374 89118 120000 89178
rect 117926 88438 120000 88498
rect 0 87758 1306 87818
rect 118202 87758 120000 87818
rect 0 87078 1490 87138
rect 0 86398 846 86458
rect 118110 86398 120000 86458
rect 117834 85718 120000 85778
rect 0 85038 754 85098
rect 117742 85038 120000 85098
rect 0 84358 1858 84418
rect 0 83678 386 83738
rect 117834 83678 120000 83738
rect 118018 82998 120000 83058
rect 0 82318 754 82378
rect 0 81638 1858 81698
rect 117190 81638 120000 81698
rect 0 80958 754 81018
rect 118110 80958 120000 81018
rect 118110 80278 120000 80338
rect 0 79598 846 79658
rect 0 78918 1582 78978
rect 118110 78918 120000 78978
rect 117834 78238 120000 78298
rect 0 77558 662 77618
rect 118110 77558 120000 77618
rect 0 76878 1858 76938
rect 0 76198 1306 76258
rect 117834 76198 120000 76258
rect 118110 75518 120000 75578
rect 0 74838 662 74898
rect 0 74158 1306 74218
rect 117834 74158 120000 74218
rect 0 73478 754 73538
rect 118110 73478 120000 73538
rect 118110 72798 120000 72858
rect 0 72118 1398 72178
rect 0 71438 1398 71498
rect 118110 71438 120000 71498
rect 117926 70758 120000 70818
rect 0 70078 1306 70138
rect 118110 70078 120000 70138
rect 0 69398 754 69458
rect 0 68718 1306 68778
rect 117834 68718 120000 68778
rect 118110 68038 120000 68098
rect 0 67358 1398 67418
rect 118110 67358 120000 67418
rect 0 66678 754 66738
rect 0 65998 1122 66058
rect 118202 65998 120000 66058
rect 117926 65318 120000 65378
rect 0 64638 1490 64698
rect 0 63958 1214 64018
rect 117926 63958 120000 64018
rect 0 63278 846 63338
rect 117926 63278 120000 63338
rect 118110 62598 120000 62658
rect 0 61918 754 61978
rect 0 61238 754 61298
rect 118110 61238 120000 61298
rect 118202 60558 120000 60618
rect 0 59878 1306 59938
rect 118110 59878 120000 59938
rect 0 59198 1306 59258
rect 0 58518 754 58578
rect 118110 58518 120000 58578
rect 117834 57838 120000 57898
rect 0 57158 1122 57218
rect 0 56478 754 56538
rect 117926 56478 120000 56538
rect 0 55798 1306 55858
rect 118110 55798 120000 55858
rect 118110 55118 120000 55178
rect 0 54438 1398 54498
rect 0 53758 1490 53818
rect 117374 53758 120000 53818
rect 117834 53078 120000 53138
rect 0 52398 846 52458
rect 117926 52398 120000 52458
rect 0 51718 386 51778
rect 0 51038 1398 51098
rect 117834 51038 120000 51098
rect 118110 50358 120000 50418
rect 0 49678 386 49738
rect 118202 49678 120000 49738
rect 0 48998 386 49058
rect 0 48318 1582 48378
rect 118110 48318 120000 48378
rect 118110 47638 120000 47698
rect 0 46958 1490 47018
rect 0 46278 386 46338
rect 118018 46278 120000 46338
rect 0 45598 1490 45658
rect 117834 45598 120000 45658
rect 117926 44918 120000 44978
rect 0 44238 1306 44298
rect 0 43558 1398 43618
rect 117742 43558 120000 43618
rect 118110 42878 120000 42938
rect 0 42198 1306 42258
rect 118110 42198 120000 42258
rect 0 41518 1306 41578
rect 0 40838 1490 40898
rect 118110 40838 120000 40898
rect 118110 40158 120000 40218
rect 0 39478 1306 39538
rect 0 38798 1122 38858
rect 118202 38798 120000 38858
rect 0 38118 386 38178
rect 117834 38118 120000 38178
rect 118110 37438 120000 37498
rect 0 36758 1306 36818
rect 0 36078 1306 36138
rect 117834 36078 120000 36138
rect 118110 35398 120000 35458
rect 0 34718 386 34778
rect 117834 34718 120000 34778
rect 0 34038 1398 34098
rect 0 33358 1122 33418
rect 118110 33358 120000 33418
rect 117834 32678 120000 32738
rect 0 31998 1306 32058
rect 118202 31998 120000 32058
rect 0 31318 1398 31378
rect 0 30638 846 30698
rect 117834 30638 120000 30698
rect 118110 29958 120000 30018
rect 0 29278 386 29338
rect 0 28598 1582 28658
rect 118110 28598 120000 28658
rect 0 27918 1122 27978
rect 118110 27918 120000 27978
rect 117834 27238 120000 27298
rect 0 26558 386 26618
rect 0 25878 1490 25938
rect 117834 25878 120000 25938
rect 117834 25198 120000 25258
rect 0 24518 1858 24578
rect 118202 24518 120000 24578
rect 0 23838 1306 23898
rect 0 23158 662 23218
rect 117926 23158 120000 23218
rect 118202 22478 120000 22538
rect 0 21798 1398 21858
rect 0 21118 1306 21178
rect 118110 21118 120000 21178
rect 0 20438 1398 20498
rect 118110 20438 120000 20498
rect 117742 19758 120000 19818
rect 0 19078 386 19138
rect 0 18398 846 18458
rect 117834 18398 120000 18458
rect 118110 17718 120000 17778
rect 0 17038 386 17098
rect 118110 17038 120000 17098
rect 0 16358 1306 16418
rect 0 15678 1582 15738
rect 118110 15678 120000 15738
rect 118110 14998 120000 15058
rect 0 14318 846 14378
rect 117834 14318 120000 14378
rect 0 13638 754 13698
rect 0 12958 1490 13018
rect 117926 12958 120000 13018
rect 118202 12278 120000 12338
rect 0 11598 754 11658
rect 0 10918 1858 10978
rect 117926 10918 120000 10978
rect 0 10238 386 10298
rect 118202 10238 120000 10298
rect 117834 9558 120000 9618
rect 0 8878 1306 8938
rect 0 8198 1490 8258
rect 118202 8198 120000 8258
rect 117834 7518 120000 7578
rect 0 6838 1582 6898
rect 118110 6838 120000 6898
rect 0 6158 754 6218
rect 0 5478 1582 5538
rect 117834 5478 120000 5538
rect 118110 4798 120000 4858
rect 0 4118 1306 4178
rect 0 3438 1306 3498
rect 117098 3438 120000 3498
rect 0 2758 754 2818
rect 117374 2758 120000 2818
rect 118018 2078 120000 2138
rect 0 1398 1122 1458
rect 0 718 2226 778
rect 116638 718 120000 778
rect 119214 38 120000 98
<< obsm3 >>
rect 1478 119638 119219 119781
rect 381 119178 119219 119638
rect 1570 118958 117846 119178
rect 381 118498 119219 118958
rect 381 118278 116190 118498
rect 381 117818 119219 118278
rect 2306 117598 119219 117818
rect 381 117138 119219 117598
rect 2858 116918 117294 117138
rect 381 116458 119219 116918
rect 926 116238 117754 116458
rect 381 115778 119219 116238
rect 381 115558 118030 115778
rect 381 115098 119219 115558
rect 1938 114878 119219 115098
rect 381 114418 119219 114878
rect 1386 114198 117754 114418
rect 381 113738 119219 114198
rect 381 113518 118030 113738
rect 381 113058 119219 113518
rect 650 112838 117754 113058
rect 381 112378 119219 112838
rect 1386 112158 119219 112378
rect 381 111698 119219 112158
rect 466 111478 118030 111698
rect 381 111018 119219 111478
rect 381 110798 117252 111018
rect 381 110338 119219 110798
rect 834 110118 119219 110338
rect 381 109658 119219 110118
rect 1386 109438 118030 109658
rect 381 108978 119219 109438
rect 1478 108758 117846 108978
rect 381 108298 119219 108758
rect 381 108078 118030 108298
rect 381 107618 119219 108078
rect 1386 107398 119219 107618
rect 381 106938 119219 107398
rect 926 106718 117754 106938
rect 381 106258 119219 106718
rect 381 106038 118030 106258
rect 381 105578 119219 106038
rect 1570 105358 117662 105578
rect 381 104898 119219 105358
rect 834 104678 119219 104898
rect 381 104218 119219 104678
rect 466 103998 118030 104218
rect 381 103538 119219 103998
rect 381 103318 117754 103538
rect 381 102858 119219 103318
rect 1570 102638 118030 102858
rect 381 102178 119219 102638
rect 742 101958 119219 102178
rect 381 101498 119219 101958
rect 1386 101278 117754 101498
rect 381 100818 119219 101278
rect 381 100598 118030 100818
rect 381 100138 119219 100598
rect 1478 99918 119219 100138
rect 381 99458 119219 99918
rect 1662 99238 118030 99458
rect 381 98778 119219 99238
rect 466 98558 118122 98778
rect 381 98098 119219 98558
rect 381 97878 117754 98098
rect 381 97418 119219 97878
rect 466 97198 119219 97418
rect 381 96738 119219 97198
rect 1570 96518 117754 96738
rect 381 96058 119219 96518
rect 381 95838 118030 96058
rect 381 95378 119219 95838
rect 1202 95158 117754 95378
rect 381 94698 119219 95158
rect 466 94478 119219 94698
rect 381 94018 119219 94478
rect 742 93798 117018 94018
rect 381 93338 119219 93798
rect 381 93118 116190 93338
rect 381 92658 119219 93118
rect 466 92438 119219 92658
rect 381 91978 119219 92438
rect 926 91758 116834 91978
rect 381 91298 119219 91758
rect 1478 91078 118030 91298
rect 381 90618 119219 91078
rect 381 90398 117754 90618
rect 381 89938 119219 90398
rect 1570 89718 119219 89938
rect 381 89258 119219 89718
rect 926 89038 117294 89258
rect 381 88578 119219 89038
rect 381 88358 117846 88578
rect 381 87898 119219 88358
rect 1386 87678 118122 87898
rect 381 87218 119219 87678
rect 1570 86998 119219 87218
rect 381 86538 119219 86998
rect 926 86318 118030 86538
rect 381 85858 119219 86318
rect 381 85638 117754 85858
rect 381 85178 119219 85638
rect 834 84958 117662 85178
rect 381 84498 119219 84958
rect 1938 84278 119219 84498
rect 381 83818 119219 84278
rect 466 83598 117754 83818
rect 381 83138 119219 83598
rect 381 82918 117938 83138
rect 381 82458 119219 82918
rect 834 82238 119219 82458
rect 381 81778 119219 82238
rect 1938 81558 117110 81778
rect 381 81098 119219 81558
rect 834 80878 118030 81098
rect 381 80418 119219 80878
rect 381 80198 118030 80418
rect 381 79738 119219 80198
rect 926 79518 119219 79738
rect 381 79058 119219 79518
rect 1662 78838 118030 79058
rect 381 78378 119219 78838
rect 381 78158 117754 78378
rect 381 77698 119219 78158
rect 742 77478 118030 77698
rect 381 77018 119219 77478
rect 1938 76798 119219 77018
rect 381 76338 119219 76798
rect 1386 76118 117754 76338
rect 381 75658 119219 76118
rect 381 75438 118030 75658
rect 381 74978 119219 75438
rect 742 74758 119219 74978
rect 381 74298 119219 74758
rect 1386 74078 117754 74298
rect 381 73618 119219 74078
rect 834 73398 118030 73618
rect 381 72938 119219 73398
rect 381 72718 118030 72938
rect 381 72258 119219 72718
rect 1478 72038 119219 72258
rect 381 71578 119219 72038
rect 1478 71358 118030 71578
rect 381 70898 119219 71358
rect 381 70678 117846 70898
rect 381 70218 119219 70678
rect 1386 69998 118030 70218
rect 381 69538 119219 69998
rect 834 69318 119219 69538
rect 381 68858 119219 69318
rect 1386 68638 117754 68858
rect 381 68178 119219 68638
rect 381 67958 118030 68178
rect 381 67498 119219 67958
rect 1478 67278 118030 67498
rect 381 66818 119219 67278
rect 834 66598 119219 66818
rect 381 66138 119219 66598
rect 1202 65918 118122 66138
rect 381 65458 119219 65918
rect 381 65238 117846 65458
rect 381 64778 119219 65238
rect 1570 64558 119219 64778
rect 381 64098 119219 64558
rect 1294 63878 117846 64098
rect 381 63418 119219 63878
rect 926 63198 117846 63418
rect 381 62738 119219 63198
rect 381 62518 118030 62738
rect 381 62058 119219 62518
rect 834 61838 119219 62058
rect 381 61378 119219 61838
rect 834 61158 118030 61378
rect 381 60698 119219 61158
rect 381 60478 118122 60698
rect 381 60018 119219 60478
rect 1386 59798 118030 60018
rect 381 59338 119219 59798
rect 1386 59118 119219 59338
rect 381 58658 119219 59118
rect 834 58438 118030 58658
rect 381 57978 119219 58438
rect 381 57758 117754 57978
rect 381 57298 119219 57758
rect 1202 57078 119219 57298
rect 381 56618 119219 57078
rect 834 56398 117846 56618
rect 381 55938 119219 56398
rect 1386 55718 118030 55938
rect 381 55258 119219 55718
rect 381 55038 118030 55258
rect 381 54578 119219 55038
rect 1478 54358 119219 54578
rect 381 53898 119219 54358
rect 1570 53678 117294 53898
rect 381 53218 119219 53678
rect 381 52998 117754 53218
rect 381 52538 119219 52998
rect 926 52318 117846 52538
rect 381 51858 119219 52318
rect 466 51638 119219 51858
rect 381 51178 119219 51638
rect 1478 50958 117754 51178
rect 381 50498 119219 50958
rect 381 50278 118030 50498
rect 381 49818 119219 50278
rect 466 49598 118122 49818
rect 381 49138 119219 49598
rect 466 48918 119219 49138
rect 381 48458 119219 48918
rect 1662 48238 118030 48458
rect 381 47778 119219 48238
rect 381 47558 118030 47778
rect 381 47098 119219 47558
rect 1570 46878 119219 47098
rect 381 46418 119219 46878
rect 466 46198 117938 46418
rect 381 45738 119219 46198
rect 1570 45518 117754 45738
rect 381 45058 119219 45518
rect 381 44838 117846 45058
rect 381 44378 119219 44838
rect 1386 44158 119219 44378
rect 381 43698 119219 44158
rect 1478 43478 117662 43698
rect 381 43018 119219 43478
rect 381 42798 118030 43018
rect 381 42338 119219 42798
rect 1386 42118 118030 42338
rect 381 41658 119219 42118
rect 1386 41438 119219 41658
rect 381 40978 119219 41438
rect 1570 40758 118030 40978
rect 381 40298 119219 40758
rect 381 40078 118030 40298
rect 381 39618 119219 40078
rect 1386 39398 119219 39618
rect 381 38938 119219 39398
rect 1202 38718 118122 38938
rect 381 38258 119219 38718
rect 466 38038 117754 38258
rect 381 37578 119219 38038
rect 381 37358 118030 37578
rect 381 36898 119219 37358
rect 1386 36678 119219 36898
rect 381 36218 119219 36678
rect 1386 35998 117754 36218
rect 381 35538 119219 35998
rect 381 35318 118030 35538
rect 381 34858 119219 35318
rect 466 34638 117754 34858
rect 381 34178 119219 34638
rect 1478 33958 119219 34178
rect 381 33498 119219 33958
rect 1202 33278 118030 33498
rect 381 32818 119219 33278
rect 381 32598 117754 32818
rect 381 32138 119219 32598
rect 1386 31918 118122 32138
rect 381 31458 119219 31918
rect 1478 31238 119219 31458
rect 381 30778 119219 31238
rect 926 30558 117754 30778
rect 381 30098 119219 30558
rect 381 29878 118030 30098
rect 381 29418 119219 29878
rect 466 29198 119219 29418
rect 381 28738 119219 29198
rect 1662 28518 118030 28738
rect 381 28058 119219 28518
rect 1202 27838 118030 28058
rect 381 27378 119219 27838
rect 381 27158 117754 27378
rect 381 26698 119219 27158
rect 466 26478 119219 26698
rect 381 26018 119219 26478
rect 1570 25798 117754 26018
rect 381 25338 119219 25798
rect 381 25118 117754 25338
rect 381 24658 119219 25118
rect 1938 24438 118122 24658
rect 381 23978 119219 24438
rect 1386 23758 119219 23978
rect 381 23298 119219 23758
rect 742 23078 117846 23298
rect 381 22618 119219 23078
rect 381 22398 118122 22618
rect 381 21938 119219 22398
rect 1478 21718 119219 21938
rect 381 21258 119219 21718
rect 1386 21038 118030 21258
rect 381 20578 119219 21038
rect 1478 20358 118030 20578
rect 381 19898 119219 20358
rect 381 19678 117662 19898
rect 381 19218 119219 19678
rect 466 18998 119219 19218
rect 381 18538 119219 18998
rect 926 18318 117754 18538
rect 381 17858 119219 18318
rect 381 17638 118030 17858
rect 381 17178 119219 17638
rect 466 16958 118030 17178
rect 381 16498 119219 16958
rect 1386 16278 119219 16498
rect 381 15818 119219 16278
rect 1662 15598 118030 15818
rect 381 15138 119219 15598
rect 381 14918 118030 15138
rect 381 14458 119219 14918
rect 926 14238 117754 14458
rect 381 13778 119219 14238
rect 834 13558 119219 13778
rect 381 13098 119219 13558
rect 1570 12878 117846 13098
rect 381 12418 119219 12878
rect 381 12198 118122 12418
rect 381 11738 119219 12198
rect 834 11518 119219 11738
rect 381 11058 119219 11518
rect 1938 10838 117846 11058
rect 381 10378 119219 10838
rect 466 10158 118122 10378
rect 381 9698 119219 10158
rect 381 9478 117754 9698
rect 381 9018 119219 9478
rect 1386 8798 119219 9018
rect 381 8338 119219 8798
rect 1570 8118 118122 8338
rect 381 7658 119219 8118
rect 381 7438 117754 7658
rect 381 6978 119219 7438
rect 1662 6758 118030 6978
rect 381 6298 119219 6758
rect 834 6078 119219 6298
rect 381 5618 119219 6078
rect 1662 5398 117754 5618
rect 381 4938 119219 5398
rect 381 4718 118030 4938
rect 381 4258 119219 4718
rect 1386 4038 119219 4258
rect 381 3578 119219 4038
rect 1386 3358 117018 3578
rect 381 2898 119219 3358
rect 834 2678 117294 2898
rect 381 2218 119219 2678
rect 381 1998 117938 2218
rect 381 1538 119219 1998
rect 1202 1318 119219 1538
rect 381 858 119219 1318
rect 2306 638 116558 858
rect 381 178 119219 638
rect 381 35 119134 178
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 1262 2262 4128 117197
rect 4608 2262 19488 117197
rect 19968 2262 34848 117197
rect 35328 2262 50208 117197
rect 50688 2262 65568 117197
rect 66048 2262 80928 117197
rect 81408 2262 96288 117197
rect 96768 2262 111648 117197
rect 112128 2262 118069 117197
<< metal5 >>
rect 1056 112572 118912 112892
rect 1056 97254 118912 97574
rect 1056 81936 118912 82256
rect 1056 66618 118912 66938
rect 1056 51300 118912 51620
rect 1056 35982 118912 36302
rect 1056 20664 118912 20984
rect 1056 5346 118912 5666
<< obsm5 >>
rect 1220 113212 117828 116780
rect 1220 97894 117828 112252
rect 1220 82576 117828 96934
rect 1220 67258 117828 81616
rect 1220 51940 117828 66298
rect 1220 36622 117828 50980
rect 1220 21304 117828 35662
rect 1220 5986 117828 20344
rect 1220 2220 117828 5026
<< labels >>
rlabel metal3 s 117332 110878 120000 110938 6 clk
port 1 nsew signal input
rlabel metal3 s 0 36758 1306 36818 6 enable
port 2 nsew signal input
rlabel metal3 s 118110 80958 120000 81018 6 finish
port 3 nsew signal output
rlabel metal3 s 0 107478 1306 107538 6 rst
port 4 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 5346 118912 5666 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 35982 118912 36302 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 66618 118912 66938 6 vccd1
port 5 nsew power bidirectional
rlabel metal5 s 1056 97254 118912 97574 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 20664 118912 20984 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 51300 118912 51620 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 81936 118912 82256 6 vssd1
port 6 nsew ground bidirectional
rlabel metal5 s 1056 112572 118912 112892 6 vssd1
port 6 nsew ground bidirectional
rlabel metal2 s 7116 117292 7144 120000 6 x_i_0[0]
port 7 nsew signal input
rlabel metal2 s 20640 117292 20668 120000 6 x_i_0[10]
port 8 nsew signal input
rlabel metal3 s 0 81638 1858 81698 6 x_i_0[11]
port 9 nsew signal input
rlabel metal3 s 118202 24518 120000 24578 6 x_i_0[12]
port 10 nsew signal input
rlabel metal3 s 118110 48318 120000 48378 6 x_i_0[13]
port 11 nsew signal input
rlabel metal3 s 118110 29958 120000 30018 6 x_i_0[14]
port 12 nsew signal input
rlabel metal3 s 118110 67358 120000 67418 6 x_i_0[15]
port 13 nsew signal input
rlabel metal2 s 22572 0 22600 2388 6 x_i_0[1]
port 14 nsew signal input
rlabel metal3 s 0 55798 1306 55858 6 x_i_0[2]
port 15 nsew signal input
rlabel metal3 s 0 84358 1858 84418 6 x_i_0[3]
port 16 nsew signal input
rlabel metal2 s 106936 0 106964 3000 6 x_i_0[4]
port 17 nsew signal input
rlabel metal3 s 117834 36078 120000 36138 6 x_i_0[5]
port 18 nsew signal input
rlabel metal3 s 0 78918 1582 78978 6 x_i_0[6]
port 19 nsew signal input
rlabel metal3 s 0 72118 1398 72178 6 x_i_0[7]
port 20 nsew signal input
rlabel metal2 s 117240 117292 117268 120000 6 x_i_0[8]
port 21 nsew signal input
rlabel metal3 s 117834 76198 120000 76258 6 x_i_0[9]
port 22 nsew signal input
rlabel metal3 s 118202 38798 120000 38858 6 x_i_1[0]
port 23 nsew signal input
rlabel metal2 s 82464 0 82492 218 6 x_i_1[10]
port 24 nsew signal input
rlabel metal2 s 21928 0 21956 2320 6 x_i_1[11]
port 25 nsew signal input
rlabel metal2 s 3252 0 3280 3000 6 x_i_1[12]
port 26 nsew signal input
rlabel metal2 s 55416 0 55444 2258 6 x_i_1[13]
port 27 nsew signal input
rlabel metal3 s 117834 18398 120000 18458 6 x_i_1[14]
port 28 nsew signal input
rlabel metal3 s 117374 53758 120000 53818 6 x_i_1[15]
port 29 nsew signal input
rlabel metal2 s 43824 0 43852 2388 6 x_i_1[1]
port 30 nsew signal input
rlabel metal3 s 0 4118 1306 4178 6 x_i_1[2]
port 31 nsew signal input
rlabel metal3 s 0 21118 1306 21178 6 x_i_1[3]
port 32 nsew signal input
rlabel metal2 s 41892 117292 41920 120000 6 x_i_1[4]
port 33 nsew signal input
rlabel metal3 s 118202 65998 120000 66058 6 x_i_1[5]
port 34 nsew signal input
rlabel metal3 s 117926 65318 120000 65378 6 x_i_1[6]
port 35 nsew signal input
rlabel metal2 s 6472 116680 6500 120000 6 x_i_1[7]
port 36 nsew signal input
rlabel metal3 s 118202 98638 120000 98698 6 x_i_1[8]
port 37 nsew signal input
rlabel metal3 s 0 44238 1306 44298 6 x_i_1[9]
port 38 nsew signal input
rlabel metal3 s 116914 91838 120000 91898 6 x_i_2[0]
port 39 nsew signal input
rlabel metal2 s 108868 117292 108896 120000 6 x_i_2[10]
port 40 nsew signal input
rlabel metal2 s 18064 0 18092 2388 6 x_i_2[11]
port 41 nsew signal input
rlabel metal2 s 112732 0 112760 2388 6 x_i_2[12]
port 42 nsew signal input
rlabel metal2 s 52196 116680 52224 120000 6 x_i_2[13]
port 43 nsew signal input
rlabel metal2 s 33520 0 33548 2388 6 x_i_2[14]
port 44 nsew signal input
rlabel metal3 s 0 119038 1490 119098 6 x_i_2[15]
port 45 nsew signal input
rlabel metal2 s 101140 0 101168 3000 6 x_i_2[1]
port 46 nsew signal input
rlabel metal2 s 39316 116680 39344 120000 6 x_i_2[2]
port 47 nsew signal input
rlabel metal3 s 0 67358 1398 67418 6 x_i_2[3]
port 48 nsew signal input
rlabel metal2 s 36096 0 36124 2320 6 x_i_2[4]
port 49 nsew signal input
rlabel metal2 s 67008 117292 67036 120000 6 x_i_2[5]
port 50 nsew signal input
rlabel metal2 s 54772 117292 54800 120000 6 x_i_2[6]
port 51 nsew signal input
rlabel metal3 s 0 15678 1582 15738 6 x_i_2[7]
port 52 nsew signal input
rlabel metal3 s 0 70078 1306 70138 6 x_i_2[8]
port 53 nsew signal input
rlabel metal2 s 77312 0 77340 2320 6 x_i_2[9]
port 54 nsew signal input
rlabel metal3 s 0 34038 1398 34098 6 x_i_3[0]
port 55 nsew signal input
rlabel metal2 s 7760 0 7788 2320 6 x_i_3[10]
port 56 nsew signal input
rlabel metal2 s 13556 116680 13584 120000 6 x_i_3[11]
port 57 nsew signal input
rlabel metal3 s 118110 55798 120000 55858 6 x_i_3[12]
port 58 nsew signal input
rlabel metal3 s 0 65998 1122 66058 6 x_i_3[13]
port 59 nsew signal input
rlabel metal2 s 100496 119870 100524 120000 6 x_i_3[14]
port 60 nsew signal input
rlabel metal3 s 0 87758 1306 87818 6 x_i_3[15]
port 61 nsew signal input
rlabel metal3 s 117926 108838 120000 108898 6 x_i_3[1]
port 62 nsew signal input
rlabel metal2 s 119816 0 119844 1300 6 x_i_3[2]
port 63 nsew signal input
rlabel metal2 s 57992 0 58020 2388 6 x_i_3[3]
port 64 nsew signal input
rlabel metal2 s 118528 117428 118556 120000 6 x_i_3[4]
port 65 nsew signal input
rlabel metal3 s 116270 93198 120000 93258 6 x_i_3[5]
port 66 nsew signal input
rlabel metal2 s 2608 119870 2636 120000 6 x_i_3[6]
port 67 nsew signal input
rlabel metal2 s 110800 0 110828 3000 6 x_i_3[7]
port 68 nsew signal input
rlabel metal2 s 56060 116884 56088 120000 6 x_i_3[8]
port 69 nsew signal input
rlabel metal3 s 0 41518 1306 41578 6 x_i_3[9]
port 70 nsew signal input
rlabel metal2 s 75380 0 75408 2258 6 x_i_4[0]
port 71 nsew signal input
rlabel metal3 s 0 71438 1398 71498 6 x_i_4[10]
port 72 nsew signal input
rlabel metal2 s 114020 117292 114048 120000 6 x_i_4[11]
port 73 nsew signal input
rlabel metal3 s 0 5478 1582 5538 6 x_i_4[12]
port 74 nsew signal input
rlabel metal2 s 74736 0 74764 2388 6 x_i_4[13]
port 75 nsew signal input
rlabel metal2 s 39960 0 39988 2320 6 x_i_4[14]
port 76 nsew signal input
rlabel metal3 s 0 38798 1122 38858 6 x_i_4[15]
port 77 nsew signal input
rlabel metal3 s 118202 12278 120000 12338 6 x_i_4[1]
port 78 nsew signal input
rlabel metal3 s 118110 14998 120000 15058 6 x_i_4[2]
port 79 nsew signal input
rlabel metal3 s 118110 58518 120000 58578 6 x_i_4[3]
port 80 nsew signal input
rlabel metal3 s 118110 109518 120000 109578 6 x_i_4[4]
port 81 nsew signal input
rlabel metal3 s 0 59198 1306 59258 6 x_i_4[5]
port 82 nsew signal input
rlabel metal2 s 41248 0 41276 2252 6 x_i_4[6]
port 83 nsew signal input
rlabel metal3 s 0 57158 1122 57218 6 x_i_4[7]
port 84 nsew signal input
rlabel metal2 s 111444 0 111472 2320 6 x_i_4[8]
port 85 nsew signal input
rlabel metal3 s 0 54438 1398 54498 6 x_i_4[9]
port 86 nsew signal input
rlabel metal3 s 117926 10918 120000 10978 6 x_i_5[0]
port 87 nsew signal input
rlabel metal3 s 118110 111558 120000 111618 6 x_i_5[10]
port 88 nsew signal input
rlabel metal2 s 38028 117292 38056 120000 6 x_i_5[11]
port 89 nsew signal input
rlabel metal2 s 90836 117292 90864 120000 6 x_i_5[12]
port 90 nsew signal input
rlabel metal2 s 94700 0 94728 1300 6 x_i_5[13]
port 91 nsew signal input
rlabel metal3 s 118110 72798 120000 72858 6 x_i_5[14]
port 92 nsew signal input
rlabel metal3 s 0 112238 1306 112298 6 x_i_5[15]
port 93 nsew signal input
rlabel metal2 s 52840 0 52868 2320 6 x_i_5[1]
port 94 nsew signal input
rlabel metal2 s 61856 117292 61884 120000 6 x_i_5[2]
port 95 nsew signal input
rlabel metal2 s 69584 0 69612 2388 6 x_i_5[3]
port 96 nsew signal input
rlabel metal3 s 0 24518 1858 24578 6 x_i_5[4]
port 97 nsew signal input
rlabel metal2 s 87616 117292 87644 120000 6 x_i_5[5]
port 98 nsew signal input
rlabel metal3 s 118110 59878 120000 59938 6 x_i_5[6]
port 99 nsew signal input
rlabel metal3 s 0 16358 1306 16418 6 x_i_5[7]
port 100 nsew signal input
rlabel metal3 s 118110 42198 120000 42258 6 x_i_5[8]
port 101 nsew signal input
rlabel metal3 s 0 101358 1306 101418 6 x_i_5[9]
port 102 nsew signal input
rlabel metal3 s 117098 3438 120000 3498 6 x_i_6[0]
port 103 nsew signal input
rlabel metal3 s 0 6838 1582 6898 6 x_i_6[10]
port 104 nsew signal input
rlabel metal3 s 0 21798 1398 21858 6 x_i_6[11]
port 105 nsew signal input
rlabel metal3 s 0 51038 1398 51098 6 x_i_6[12]
port 106 nsew signal input
rlabel metal2 s 74092 117292 74120 120000 6 x_i_6[13]
port 107 nsew signal input
rlabel metal2 s 19352 117292 19380 120000 6 x_i_6[14]
port 108 nsew signal input
rlabel metal3 s 118202 22478 120000 22538 6 x_i_6[15]
port 109 nsew signal input
rlabel metal2 s 61212 0 61240 2388 6 x_i_6[1]
port 110 nsew signal input
rlabel metal3 s 0 36078 1306 36138 6 x_i_6[2]
port 111 nsew signal input
rlabel metal2 s 16132 117292 16160 120000 6 x_i_6[3]
port 112 nsew signal input
rlabel metal3 s 0 42198 1306 42258 6 x_i_6[4]
port 113 nsew signal input
rlabel metal2 s 49620 116680 49648 120000 6 x_i_6[5]
port 114 nsew signal input
rlabel metal2 s 29656 0 29684 2320 6 x_i_6[6]
port 115 nsew signal input
rlabel metal3 s 118110 61238 120000 61298 6 x_i_6[7]
port 116 nsew signal input
rlabel metal2 s 119172 115116 119200 120000 6 x_i_6[8]
port 117 nsew signal input
rlabel metal2 s 107580 116884 107608 120000 6 x_i_6[9]
port 118 nsew signal input
rlabel metal3 s 118110 40158 120000 40218 6 x_i_7[0]
port 119 nsew signal input
rlabel metal2 s 68296 0 68324 1300 6 x_i_7[10]
port 120 nsew signal input
rlabel metal3 s 118110 20438 120000 20498 6 x_i_7[11]
port 121 nsew signal input
rlabel metal2 s 97920 117360 97948 120000 6 x_i_7[12]
port 122 nsew signal input
rlabel metal2 s 113376 116680 113404 120000 6 x_i_7[13]
port 123 nsew signal input
rlabel metal3 s 0 76198 1306 76258 6 x_i_7[14]
port 124 nsew signal input
rlabel metal3 s 0 43558 1398 43618 6 x_i_7[15]
port 125 nsew signal input
rlabel metal2 s 65720 0 65748 218 6 x_i_7[1]
port 126 nsew signal input
rlabel metal3 s 118202 10238 120000 10298 6 x_i_7[2]
port 127 nsew signal input
rlabel metal2 s 16776 117292 16804 120000 6 x_i_7[3]
port 128 nsew signal input
rlabel metal3 s 118202 87758 120000 87818 6 x_i_7[4]
port 129 nsew signal input
rlabel metal2 s 17420 0 17448 2320 6 x_i_7[5]
port 130 nsew signal input
rlabel metal2 s 44468 117292 44496 120000 6 x_i_7[6]
port 131 nsew signal input
rlabel metal2 s 63144 117360 63172 120000 6 x_i_7[7]
port 132 nsew signal input
rlabel metal3 s 0 114278 1306 114338 6 x_i_7[8]
port 133 nsew signal input
rlabel metal3 s 0 31998 1306 32058 6 x_i_7[9]
port 134 nsew signal input
rlabel metal2 s 106292 117292 106320 120000 6 x_r_0[0]
port 135 nsew signal input
rlabel metal2 s 91480 0 91508 1300 6 x_r_0[10]
port 136 nsew signal input
rlabel metal2 s 47044 0 47072 2388 6 x_r_0[11]
port 137 nsew signal input
rlabel metal2 s 68940 117292 68968 120000 6 x_r_0[12]
port 138 nsew signal input
rlabel metal3 s 116638 718 120000 778 6 x_r_0[13]
port 139 nsew signal input
rlabel metal3 s 0 76878 1858 76938 6 x_r_0[14]
port 140 nsew signal input
rlabel metal2 s 36096 117292 36124 120000 6 x_r_0[15]
port 141 nsew signal input
rlabel metal3 s 117926 56478 120000 56538 6 x_r_0[1]
port 142 nsew signal input
rlabel metal3 s 0 99318 1582 99378 6 x_r_0[2]
port 143 nsew signal input
rlabel metal3 s 0 74158 1306 74218 6 x_r_0[3]
port 144 nsew signal input
rlabel metal2 s 34164 0 34192 218 6 x_r_0[4]
port 145 nsew signal input
rlabel metal2 s 41892 0 41920 2796 6 x_r_0[5]
port 146 nsew signal input
rlabel metal2 s 22572 116680 22600 120000 6 x_r_0[6]
port 147 nsew signal input
rlabel metal3 s 0 28598 1582 28658 6 x_r_0[7]
port 148 nsew signal input
rlabel metal2 s 113376 0 113404 2320 6 x_r_0[8]
port 149 nsew signal input
rlabel metal2 s 117240 0 117268 3408 6 x_r_0[9]
port 150 nsew signal input
rlabel metal2 s 72804 0 72832 218 6 x_r_1[0]
port 151 nsew signal input
rlabel metal3 s 118110 47638 120000 47698 6 x_r_1[10]
port 152 nsew signal input
rlabel metal2 s 68296 117292 68324 120000 6 x_r_1[11]
port 153 nsew signal input
rlabel metal2 s 12268 0 12296 2388 6 x_r_1[12]
port 154 nsew signal input
rlabel metal3 s 0 27918 1122 27978 6 x_r_1[13]
port 155 nsew signal input
rlabel metal3 s 118202 60558 120000 60618 6 x_r_1[14]
port 156 nsew signal input
rlabel metal2 s 34808 0 34836 2320 6 x_r_1[15]
port 157 nsew signal input
rlabel metal3 s 117926 63958 120000 64018 6 x_r_1[1]
port 158 nsew signal input
rlabel metal2 s 51552 117292 51580 120000 6 x_r_1[2]
port 159 nsew signal input
rlabel metal2 s 52840 117292 52868 120000 6 x_r_1[3]
port 160 nsew signal input
rlabel metal2 s 65720 117292 65748 120000 6 x_r_1[4]
port 161 nsew signal input
rlabel metal2 s 85040 117292 85068 120000 6 x_r_1[5]
port 162 nsew signal input
rlabel metal3 s 0 20438 1398 20498 6 x_r_1[6]
port 163 nsew signal input
rlabel metal2 s 93412 0 93440 3000 6 x_r_1[7]
port 164 nsew signal input
rlabel metal2 s 58636 117292 58664 120000 6 x_r_1[8]
port 165 nsew signal input
rlabel metal3 s 117926 44918 120000 44978 6 x_r_1[9]
port 166 nsew signal input
rlabel metal3 s 117926 52398 120000 52458 6 x_r_2[0]
port 167 nsew signal input
rlabel metal2 s 83108 116680 83136 120000 6 x_r_2[10]
port 168 nsew signal input
rlabel metal2 s 86328 116680 86356 120000 6 x_r_2[11]
port 169 nsew signal input
rlabel metal3 s 117926 70758 120000 70818 6 x_r_2[12]
port 170 nsew signal input
rlabel metal2 s 99208 119870 99236 120000 6 x_r_2[13]
port 171 nsew signal input
rlabel metal2 s 16776 0 16804 2388 6 x_r_2[14]
port 172 nsew signal input
rlabel metal2 s 110156 0 110184 2320 6 x_r_2[15]
port 173 nsew signal input
rlabel metal2 s 50908 0 50936 3000 6 x_r_2[1]
port 174 nsew signal input
rlabel metal2 s 101784 0 101812 2320 6 x_r_2[2]
port 175 nsew signal input
rlabel metal2 s 32876 117292 32904 120000 6 x_r_2[3]
port 176 nsew signal input
rlabel metal2 s 29656 116680 29684 120000 6 x_r_2[4]
port 177 nsew signal input
rlabel metal3 s 117834 25198 120000 25258 6 x_r_2[5]
port 178 nsew signal input
rlabel metal2 s 101784 117292 101812 120000 6 x_r_2[6]
port 179 nsew signal input
rlabel metal3 s 0 39478 1306 39538 6 x_r_2[7]
port 180 nsew signal input
rlabel metal2 s 119816 117360 119844 120000 6 x_r_2[8]
port 181 nsew signal input
rlabel metal2 s 108868 0 108896 218 6 x_r_2[9]
port 182 nsew signal input
rlabel metal3 s 117834 30638 120000 30698 6 x_r_3[0]
port 183 nsew signal input
rlabel metal2 s 103072 116884 103100 120000 6 x_r_3[10]
port 184 nsew signal input
rlabel metal2 s 1320 119870 1348 120000 6 x_r_3[11]
port 185 nsew signal input
rlabel metal3 s 0 109518 1306 109578 6 x_r_3[12]
port 186 nsew signal input
rlabel metal2 s 42536 116884 42564 120000 6 x_r_3[13]
port 187 nsew signal input
rlabel metal3 s 118202 49678 120000 49738 6 x_r_3[14]
port 188 nsew signal input
rlabel metal3 s 117926 12958 120000 13018 6 x_r_3[15]
port 189 nsew signal input
rlabel metal2 s 84396 0 84424 2320 6 x_r_3[1]
port 190 nsew signal input
rlabel metal2 s 99852 117292 99880 120000 6 x_r_3[2]
port 191 nsew signal input
rlabel metal3 s 0 33358 1122 33418 6 x_r_3[3]
port 192 nsew signal input
rlabel metal2 s 45112 117292 45140 120000 6 x_r_3[4]
port 193 nsew signal input
rlabel metal3 s 118110 80278 120000 80338 6 x_r_3[5]
port 194 nsew signal input
rlabel metal2 s 23216 117292 23244 120000 6 x_r_3[6]
port 195 nsew signal input
rlabel metal3 s 0 99998 1398 100058 6 x_r_3[7]
port 196 nsew signal input
rlabel metal3 s 118110 62598 120000 62658 6 x_r_3[8]
port 197 nsew signal input
rlabel metal3 s 117834 90478 120000 90538 6 x_r_3[9]
port 198 nsew signal input
rlabel metal2 s 90192 117292 90220 120000 6 x_r_4[0]
port 199 nsew signal input
rlabel metal3 s 0 63958 1214 64018 6 x_r_4[10]
port 200 nsew signal input
rlabel metal2 s 88904 0 88932 1300 6 x_r_4[11]
port 201 nsew signal input
rlabel metal2 s 75380 117292 75408 120000 6 x_r_4[12]
port 202 nsew signal input
rlabel metal3 s 0 59878 1306 59938 6 x_r_4[13]
port 203 nsew signal input
rlabel metal2 s 46400 116884 46428 120000 6 x_r_4[14]
port 204 nsew signal input
rlabel metal3 s 117926 23158 120000 23218 6 x_r_4[15]
port 205 nsew signal input
rlabel metal3 s 0 108838 1398 108898 6 x_r_4[1]
port 206 nsew signal input
rlabel metal2 s 43180 117292 43208 120000 6 x_r_4[2]
port 207 nsew signal input
rlabel metal3 s 117190 81638 120000 81698 6 x_r_4[3]
port 208 nsew signal input
rlabel metal2 s 72160 0 72188 2252 6 x_r_4[4]
port 209 nsew signal input
rlabel metal2 s 116596 117292 116624 120000 6 x_r_4[5]
port 210 nsew signal input
rlabel metal3 s 117926 63278 120000 63338 6 x_r_4[6]
port 211 nsew signal input
rlabel metal2 s 115952 0 115980 2524 6 x_r_4[7]
port 212 nsew signal input
rlabel metal2 s 86972 0 87000 2320 6 x_r_4[8]
port 213 nsew signal input
rlabel metal2 s 104360 117292 104388 120000 6 x_r_4[9]
port 214 nsew signal input
rlabel metal3 s 118202 31998 120000 32058 6 x_r_5[0]
port 215 nsew signal input
rlabel metal2 s 39960 117360 39988 120000 6 x_r_5[10]
port 216 nsew signal input
rlabel metal3 s 0 10918 1858 10978 6 x_r_5[11]
port 217 nsew signal input
rlabel metal2 s 44468 0 44496 2320 6 x_r_5[12]
port 218 nsew signal input
rlabel metal3 s 117926 88438 120000 88498 6 x_r_5[13]
port 219 nsew signal input
rlabel metal2 s 9048 117292 9076 120000 6 x_r_5[14]
port 220 nsew signal input
rlabel metal2 s 14844 0 14872 2388 6 x_r_5[15]
port 221 nsew signal input
rlabel metal2 s 59924 117292 59952 120000 6 x_r_5[1]
port 222 nsew signal input
rlabel metal2 s 114020 0 114048 1300 6 x_r_5[2]
port 223 nsew signal input
rlabel metal2 s 46400 0 46428 2796 6 x_r_5[3]
port 224 nsew signal input
rlabel metal3 s 0 31318 1398 31378 6 x_r_5[4]
port 225 nsew signal input
rlabel metal3 s 0 114958 1858 115018 6 x_r_5[5]
port 226 nsew signal input
rlabel metal2 s 87616 0 87644 2388 6 x_r_5[6]
port 227 nsew signal input
rlabel metal2 s 1964 119870 1992 120000 6 x_r_5[7]
port 228 nsew signal input
rlabel metal3 s 0 23838 1306 23898 6 x_r_5[8]
port 229 nsew signal input
rlabel metal2 s 29012 0 29040 3000 6 x_r_5[9]
port 230 nsew signal input
rlabel metal3 s 118110 17038 120000 17098 6 x_r_6[0]
port 231 nsew signal input
rlabel metal3 s 0 48318 1582 48378 6 x_r_6[10]
port 232 nsew signal input
rlabel metal2 s 110156 117292 110184 120000 6 x_r_6[11]
port 233 nsew signal input
rlabel metal2 s 64432 116884 64460 120000 6 x_r_6[12]
port 234 nsew signal input
rlabel metal2 s 27724 117292 27752 120000 6 x_r_6[13]
port 235 nsew signal input
rlabel metal2 s 92124 117292 92152 120000 6 x_r_6[14]
port 236 nsew signal input
rlabel metal3 s 0 68718 1306 68778 6 x_r_6[15]
port 237 nsew signal input
rlabel metal2 s 10336 0 10364 2388 6 x_r_6[1]
port 238 nsew signal input
rlabel metal3 s 0 3438 1306 3498 6 x_r_6[2]
port 239 nsew signal input
rlabel metal2 s 104360 0 104388 2320 6 x_r_6[3]
port 240 nsew signal input
rlabel metal3 s 0 8878 1306 8938 6 x_r_6[4]
port 241 nsew signal input
rlabel metal3 s 118202 8198 120000 8258 6 x_r_6[5]
port 242 nsew signal input
rlabel metal3 s 117834 106798 120000 106858 6 x_r_6[6]
port 243 nsew signal input
rlabel metal2 s 59280 117292 59308 120000 6 x_r_6[7]
port 244 nsew signal input
rlabel metal3 s 118110 106118 120000 106178 6 x_r_6[8]
port 245 nsew signal input
rlabel metal2 s 60568 0 60596 2320 6 x_r_6[9]
port 246 nsew signal input
rlabel metal3 s 0 95238 1122 95298 6 x_r_7[0]
port 247 nsew signal input
rlabel metal2 s 65076 0 65104 2320 6 x_r_7[10]
port 248 nsew signal input
rlabel metal3 s 118110 35398 120000 35458 6 x_r_7[11]
port 249 nsew signal input
rlabel metal2 s 15488 116680 15516 120000 6 x_r_7[12]
port 250 nsew signal input
rlabel metal3 s 118110 33358 120000 33418 6 x_r_7[13]
port 251 nsew signal input
rlabel metal2 s 54128 0 54156 2388 6 x_r_7[14]
port 252 nsew signal input
rlabel metal2 s 53484 0 53512 218 6 x_r_7[15]
port 253 nsew signal input
rlabel metal2 s 35452 116680 35480 120000 6 x_r_7[1]
port 254 nsew signal input
rlabel metal2 s 94700 117292 94728 120000 6 x_r_7[2]
port 255 nsew signal input
rlabel metal3 s 0 91158 1398 91218 6 x_r_7[3]
port 256 nsew signal input
rlabel metal2 s 13556 0 13584 2320 6 x_r_7[4]
port 257 nsew signal input
rlabel metal2 s 81820 0 81848 490 6 x_r_7[5]
port 258 nsew signal input
rlabel metal2 s 66364 117292 66392 120000 6 x_r_7[6]
port 259 nsew signal input
rlabel metal3 s 118110 40838 120000 40898 6 x_r_7[7]
port 260 nsew signal input
rlabel metal2 s 57348 117292 57376 120000 6 x_r_7[8]
port 261 nsew signal input
rlabel metal2 s 23860 116680 23888 120000 6 x_r_7[9]
port 262 nsew signal input
rlabel metal2 s 50264 0 50292 1170 6 y_i_0[0]
port 263 nsew signal output
rlabel metal2 s 111444 117156 111472 120000 6 y_i_0[10]
port 264 nsew signal output
rlabel metal3 s 0 69398 754 69458 6 y_i_0[11]
port 265 nsew signal output
rlabel metal3 s 117834 103398 120000 103458 6 y_i_0[12]
port 266 nsew signal output
rlabel metal2 s 105004 117156 105032 120000 6 y_i_0[13]
port 267 nsew signal output
rlabel metal2 s 77956 0 77984 348 6 y_i_0[14]
port 268 nsew signal output
rlabel metal2 s 62500 0 62528 2252 6 y_i_0[15]
port 269 nsew signal output
rlabel metal2 s 27724 0 27752 2252 6 y_i_0[16]
port 270 nsew signal output
rlabel metal3 s 0 63278 846 63338 6 y_i_0[1]
port 271 nsew signal output
rlabel metal2 s 51552 0 51580 2252 6 y_i_0[2]
port 272 nsew signal output
rlabel metal2 s 4540 117156 4568 120000 6 y_i_0[3]
port 273 nsew signal output
rlabel metal3 s 0 94558 386 94618 6 y_i_0[4]
port 274 nsew signal output
rlabel metal3 s 117834 7518 120000 7578 6 y_i_0[5]
port 275 nsew signal output
rlabel metal3 s 118018 2078 120000 2138 6 y_i_0[6]
port 276 nsew signal output
rlabel metal2 s 70872 117156 70900 120000 6 y_i_0[7]
port 277 nsew signal output
rlabel metal2 s 676 0 704 1300 6 y_i_0[8]
port 278 nsew signal output
rlabel metal2 s 73448 0 73476 2252 6 y_i_0[9]
port 279 nsew signal output
rlabel metal3 s 0 93878 662 93938 6 y_i_1[0]
port 280 nsew signal output
rlabel metal2 s 40604 117156 40632 120000 6 y_i_1[10]
port 281 nsew signal output
rlabel metal3 s 0 46958 1490 47018 6 y_i_1[11]
port 282 nsew signal output
rlabel metal3 s 0 25878 1490 25938 6 y_i_1[12]
port 283 nsew signal output
rlabel metal2 s 105648 0 105676 280 6 y_i_1[13]
port 284 nsew signal output
rlabel metal3 s 0 49678 386 49738 6 y_i_1[14]
port 285 nsew signal output
rlabel metal2 s 76024 117156 76052 120000 6 y_i_1[15]
port 286 nsew signal output
rlabel metal3 s 0 102718 1490 102778 6 y_i_1[16]
port 287 nsew signal output
rlabel metal2 s 9692 116884 9720 120000 6 y_i_1[1]
port 288 nsew signal output
rlabel metal2 s 69584 117156 69612 120000 6 y_i_1[2]
port 289 nsew signal output
rlabel metal3 s 0 2758 754 2818 6 y_i_1[3]
port 290 nsew signal output
rlabel metal2 s 89548 0 89576 1170 6 y_i_1[4]
port 291 nsew signal output
rlabel metal3 s 118110 113598 120000 113658 6 y_i_1[5]
port 292 nsew signal output
rlabel metal2 s 32232 116884 32260 120000 6 y_i_1[6]
port 293 nsew signal output
rlabel metal3 s 118110 91158 120000 91218 6 y_i_1[7]
port 294 nsew signal output
rlabel metal3 s 0 48998 386 49058 6 y_i_1[8]
port 295 nsew signal output
rlabel metal3 s 117742 19758 120000 19818 6 y_i_1[9]
port 296 nsew signal output
rlabel metal3 s 0 64638 1490 64698 6 y_i_2[0]
port 297 nsew signal output
rlabel metal2 s 48976 117156 49004 120000 6 y_i_2[10]
port 298 nsew signal output
rlabel metal2 s 108224 0 108252 1164 6 y_i_2[11]
port 299 nsew signal output
rlabel metal3 s 0 74838 662 74898 6 y_i_2[12]
port 300 nsew signal output
rlabel metal2 s 5828 117156 5856 120000 6 y_i_2[13]
port 301 nsew signal output
rlabel metal3 s 117834 96598 120000 96658 6 y_i_2[14]
port 302 nsew signal output
rlabel metal3 s 0 104078 386 104138 6 y_i_2[15]
port 303 nsew signal output
rlabel metal3 s 117374 116998 120000 117058 6 y_i_2[16]
port 304 nsew signal output
rlabel metal2 s 27080 0 27108 2252 6 y_i_2[1]
port 305 nsew signal output
rlabel metal3 s 0 96598 1490 96658 6 y_i_2[2]
port 306 nsew signal output
rlabel metal2 s 80532 117156 80560 120000 6 y_i_2[3]
port 307 nsew signal output
rlabel metal3 s 118110 102718 120000 102778 6 y_i_2[4]
port 308 nsew signal output
rlabel metal3 s 118110 50358 120000 50418 6 y_i_2[5]
port 309 nsew signal output
rlabel metal3 s 0 56478 754 56538 6 y_i_2[6]
port 310 nsew signal output
rlabel metal2 s 18064 117156 18092 120000 6 y_i_2[7]
port 311 nsew signal output
rlabel metal2 s 43180 0 43208 2796 6 y_i_2[8]
port 312 nsew signal output
rlabel metal3 s 118110 73478 120000 73538 6 y_i_2[9]
port 313 nsew signal output
rlabel metal3 s 0 89118 846 89178 6 y_i_3[0]
port 314 nsew signal output
rlabel metal3 s 118018 46278 120000 46338 6 y_i_3[10]
port 315 nsew signal output
rlabel metal2 s 20640 0 20668 1170 6 y_i_3[11]
port 316 nsew signal output
rlabel metal2 s 63788 117156 63816 120000 6 y_i_3[12]
port 317 nsew signal output
rlabel metal2 s 63144 0 63172 218 6 y_i_3[13]
port 318 nsew signal output
rlabel metal2 s 56060 0 56088 2796 6 y_i_3[14]
port 319 nsew signal output
rlabel metal3 s 0 116318 846 116378 6 y_i_3[15]
port 320 nsew signal output
rlabel metal3 s 0 14318 846 14378 6 y_i_3[16]
port 321 nsew signal output
rlabel metal2 s 115308 0 115336 1028 6 y_i_3[1]
port 322 nsew signal output
rlabel metal2 s 50264 118510 50292 120000 6 y_i_3[2]
port 323 nsew signal output
rlabel metal3 s 0 91838 846 91898 6 y_i_3[3]
port 324 nsew signal output
rlabel metal2 s 39316 0 39344 2796 6 y_i_3[4]
port 325 nsew signal output
rlabel metal2 s 95344 117156 95372 120000 6 y_i_3[5]
port 326 nsew signal output
rlabel metal3 s 118018 82998 120000 83058 6 y_i_3[6]
port 327 nsew signal output
rlabel metal2 s 30300 117428 30328 120000 6 y_i_3[7]
port 328 nsew signal output
rlabel metal3 s 117742 43558 120000 43618 6 y_i_3[8]
port 329 nsew signal output
rlabel metal2 s 90192 0 90220 2796 6 y_i_3[9]
port 330 nsew signal output
rlabel metal3 s 118110 17718 120000 17778 6 y_i_4[0]
port 331 nsew signal output
rlabel metal3 s 118110 68038 120000 68098 6 y_i_4[10]
port 332 nsew signal output
rlabel metal3 s 0 111558 386 111618 6 y_i_4[11]
port 333 nsew signal output
rlabel metal3 s 0 19078 386 19138 6 y_i_4[12]
port 334 nsew signal output
rlabel metal2 s 58636 0 58664 2252 6 y_i_4[13]
port 335 nsew signal output
rlabel metal2 s 31588 0 31616 2252 6 y_i_4[14]
port 336 nsew signal output
rlabel metal3 s 117834 9558 120000 9618 6 y_i_4[15]
port 337 nsew signal output
rlabel metal2 s 6472 0 6500 2252 6 y_i_4[16]
port 338 nsew signal output
rlabel metal3 s 0 104758 754 104818 6 y_i_4[1]
port 339 nsew signal output
rlabel metal3 s 0 80958 754 81018 6 y_i_4[2]
port 340 nsew signal output
rlabel metal2 s 37384 117156 37412 120000 6 y_i_4[3]
port 341 nsew signal output
rlabel metal3 s 0 66678 754 66738 6 y_i_4[4]
port 342 nsew signal output
rlabel metal3 s 0 92518 386 92578 6 y_i_4[5]
port 343 nsew signal output
rlabel metal3 s 0 98638 386 98698 6 y_i_4[6]
port 344 nsew signal output
rlabel metal2 s 76668 0 76696 2252 6 y_i_4[7]
port 345 nsew signal output
rlabel metal3 s 117926 119038 120000 119098 6 y_i_4[8]
port 346 nsew signal output
rlabel metal3 s 0 106798 846 106858 6 y_i_4[9]
port 347 nsew signal output
rlabel metal3 s 117834 53078 120000 53138 6 y_i_5[0]
port 348 nsew signal output
rlabel metal3 s 117742 105438 120000 105498 6 y_i_5[10]
port 349 nsew signal output
rlabel metal3 s 116270 118358 120000 118418 6 y_i_5[11]
port 350 nsew signal output
rlabel metal2 s 93412 117156 93440 120000 6 y_i_5[12]
port 351 nsew signal output
rlabel metal3 s 118110 104078 120000 104138 6 y_i_5[13]
port 352 nsew signal output
rlabel metal2 s 26436 117156 26464 120000 6 y_i_5[14]
port 353 nsew signal output
rlabel metal2 s 36740 0 36768 2796 6 y_i_5[15]
port 354 nsew signal output
rlabel metal2 s 33520 117156 33548 120000 6 y_i_5[16]
port 355 nsew signal output
rlabel metal3 s 118110 27918 120000 27978 6 y_i_5[1]
port 356 nsew signal output
rlabel metal3 s 0 73478 754 73538 6 y_i_5[2]
port 357 nsew signal output
rlabel metal2 s 28368 117156 28396 120000 6 y_i_5[3]
port 358 nsew signal output
rlabel metal2 s 86328 0 86356 2796 6 y_i_5[4]
port 359 nsew signal output
rlabel metal3 s 117742 85038 120000 85098 6 y_i_5[5]
port 360 nsew signal output
rlabel metal3 s 118110 70078 120000 70138 6 y_i_5[6]
port 361 nsew signal output
rlabel metal3 s 117834 116318 120000 116378 6 y_i_5[7]
port 362 nsew signal output
rlabel metal3 s 118110 95918 120000 95978 6 y_i_5[8]
port 363 nsew signal output
rlabel metal2 s 103072 0 103100 2252 6 y_i_5[9]
port 364 nsew signal output
rlabel metal3 s 117834 97958 120000 98018 6 y_i_6[0]
port 365 nsew signal output
rlabel metal3 s 0 119718 1398 119778 6 y_i_6[10]
port 366 nsew signal output
rlabel metal2 s 118528 0 118556 3884 6 y_i_6[11]
port 367 nsew signal output
rlabel metal2 s 19996 0 20024 2252 6 y_i_6[12]
port 368 nsew signal output
rlabel metal2 s 30300 0 30328 1170 6 y_i_6[13]
port 369 nsew signal output
rlabel metal2 s 106292 0 106320 2524 6 y_i_6[14]
port 370 nsew signal output
rlabel metal3 s 117834 25878 120000 25938 6 y_i_6[15]
port 371 nsew signal output
rlabel metal3 s 118110 86398 120000 86458 6 y_i_6[16]
port 372 nsew signal output
rlabel metal2 s 76668 117156 76696 120000 6 y_i_6[1]
port 373 nsew signal output
rlabel metal2 s 71516 117428 71544 120000 6 y_i_6[2]
port 374 nsew signal output
rlabel metal2 s 54128 117156 54156 120000 6 y_i_6[3]
port 375 nsew signal output
rlabel metal3 s 0 46278 386 46338 6 y_i_6[4]
port 376 nsew signal output
rlabel metal3 s 0 97278 386 97338 6 y_i_6[5]
port 377 nsew signal output
rlabel metal3 s 0 110198 754 110258 6 y_i_6[6]
port 378 nsew signal output
rlabel metal2 s 47044 117156 47072 120000 6 y_i_6[7]
port 379 nsew signal output
rlabel metal2 s 23216 0 23244 2796 6 y_i_6[8]
port 380 nsew signal output
rlabel metal3 s 117834 85718 120000 85778 6 y_i_6[9]
port 381 nsew signal output
rlabel metal2 s 96632 117156 96660 120000 6 y_i_7[0]
port 382 nsew signal output
rlabel metal3 s 0 38118 386 38178 6 y_i_7[10]
port 383 nsew signal output
rlabel metal2 s 109512 117156 109540 120000 6 y_i_7[11]
port 384 nsew signal output
rlabel metal2 s 114664 117156 114692 120000 6 y_i_7[12]
port 385 nsew signal output
rlabel metal2 s 115952 117156 115980 120000 6 y_i_7[13]
port 386 nsew signal output
rlabel metal2 s 67008 0 67036 2252 6 y_i_7[14]
port 387 nsew signal output
rlabel metal3 s 0 6158 754 6218 6 y_i_7[15]
port 388 nsew signal output
rlabel metal2 s 3896 0 3924 2252 6 y_i_7[16]
port 389 nsew signal output
rlabel metal2 s 1320 0 1348 1170 6 y_i_7[1]
port 390 nsew signal output
rlabel metal3 s 0 82318 754 82378 6 y_i_7[2]
port 391 nsew signal output
rlabel metal3 s 0 79598 846 79658 6 y_i_7[3]
port 392 nsew signal output
rlabel metal3 s 118110 15678 120000 15738 6 y_i_7[4]
port 393 nsew signal output
rlabel metal2 s 88260 117428 88288 120000 6 y_i_7[5]
port 394 nsew signal output
rlabel metal3 s 117834 27238 120000 27298 6 y_i_7[6]
port 395 nsew signal output
rlabel metal2 s 12912 117156 12940 120000 6 y_i_7[7]
port 396 nsew signal output
rlabel metal3 s 0 61238 754 61298 6 y_i_7[8]
port 397 nsew signal output
rlabel metal2 s 25148 0 25176 2252 6 y_i_7[9]
port 398 nsew signal output
rlabel metal2 s 56704 0 56732 2252 6 y_r_0[0]
port 399 nsew signal output
rlabel metal2 s 73448 116884 73476 120000 6 y_r_0[10]
port 400 nsew signal output
rlabel metal2 s 103716 0 103744 2252 6 y_r_0[11]
port 401 nsew signal output
rlabel metal2 s 48976 0 49004 2252 6 y_r_0[12]
port 402 nsew signal output
rlabel metal2 s 96632 0 96660 2252 6 y_r_0[13]
port 403 nsew signal output
rlabel metal3 s 118110 75518 120000 75578 6 y_r_0[14]
port 404 nsew signal output
rlabel metal3 s 118110 99318 120000 99378 6 y_r_0[15]
port 405 nsew signal output
rlabel metal2 s 99208 0 99236 1170 6 y_r_0[16]
port 406 nsew signal output
rlabel metal2 s 10980 117428 11008 120000 6 y_r_0[1]
port 407 nsew signal output
rlabel metal3 s 118110 6838 120000 6898 6 y_r_0[2]
port 408 nsew signal output
rlabel metal3 s 0 89798 1490 89858 6 y_r_0[3]
port 409 nsew signal output
rlabel metal2 s 56704 117156 56732 120000 6 y_r_0[4]
port 410 nsew signal output
rlabel metal3 s 0 45598 1490 45658 6 y_r_0[5]
port 411 nsew signal output
rlabel metal2 s 97276 0 97304 2252 6 y_r_0[6]
port 412 nsew signal output
rlabel metal3 s 0 23158 662 23218 6 y_r_0[7]
port 413 nsew signal output
rlabel metal3 s 118110 21118 120000 21178 6 y_r_0[8]
port 414 nsew signal output
rlabel metal2 s 47688 117156 47716 120000 6 y_r_0[9]
port 415 nsew signal output
rlabel metal2 s 117884 0 117912 2796 6 y_r_1[0]
port 416 nsew signal output
rlabel metal2 s 3896 117156 3924 120000 6 y_r_1[10]
port 417 nsew signal output
rlabel metal2 s 15488 0 15516 2252 6 y_r_1[11]
port 418 nsew signal output
rlabel metal3 s 117834 74158 120000 74218 6 y_r_1[12]
port 419 nsew signal output
rlabel metal3 s 0 10238 386 10298 6 y_r_1[13]
port 420 nsew signal output
rlabel metal3 s 117834 95238 120000 95298 6 y_r_1[14]
port 421 nsew signal output
rlabel metal2 s 32232 0 32260 2252 6 y_r_1[15]
port 422 nsew signal output
rlabel metal3 s 0 86398 846 86458 6 y_r_1[16]
port 423 nsew signal output
rlabel metal2 s 11624 117156 11652 120000 6 y_r_1[1]
port 424 nsew signal output
rlabel metal2 s 83752 117156 83780 120000 6 y_r_1[2]
port 425 nsew signal output
rlabel metal3 s 118110 108158 120000 108218 6 y_r_1[3]
port 426 nsew signal output
rlabel metal2 s 8404 117156 8432 120000 6 y_r_1[4]
port 427 nsew signal output
rlabel metal2 s 18708 117156 18736 120000 6 y_r_1[5]
port 428 nsew signal output
rlabel metal3 s 118110 28598 120000 28658 6 y_r_1[6]
port 429 nsew signal output
rlabel metal2 s 32 115796 60 120000 6 y_r_1[7]
port 430 nsew signal output
rlabel metal3 s 117834 51038 120000 51098 6 y_r_1[8]
port 431 nsew signal output
rlabel metal3 s 0 85038 754 85098 6 y_r_1[9]
port 432 nsew signal output
rlabel metal3 s 0 17038 386 17098 6 y_r_2[0]
port 433 nsew signal output
rlabel metal3 s 0 105438 1490 105498 6 y_r_2[10]
port 434 nsew signal output
rlabel metal2 s 10980 0 11008 1170 6 y_r_2[11]
port 435 nsew signal output
rlabel metal3 s 0 61918 754 61978 6 y_r_2[12]
port 436 nsew signal output
rlabel metal3 s 117834 101358 120000 101418 6 y_r_2[13]
port 437 nsew signal output
rlabel metal3 s 0 12958 1490 13018 6 y_r_2[14]
port 438 nsew signal output
rlabel metal2 s 79244 0 79272 1164 6 y_r_2[15]
port 439 nsew signal output
rlabel metal3 s 117834 83678 120000 83738 6 y_r_2[16]
port 440 nsew signal output
rlabel metal3 s 117834 45598 120000 45658 6 y_r_2[1]
port 441 nsew signal output
rlabel metal3 s 119214 38 120000 98 6 y_r_2[2]
port 442 nsew signal output
rlabel metal3 s 0 18398 846 18458 6 y_r_2[3]
port 443 nsew signal output
rlabel metal2 s 97276 117156 97304 120000 6 y_r_2[4]
port 444 nsew signal output
rlabel metal3 s 0 51718 386 51778 6 y_r_2[5]
port 445 nsew signal output
rlabel metal2 s 100496 0 100524 218 6 y_r_2[6]
port 446 nsew signal output
rlabel metal3 s 117834 34718 120000 34778 6 y_r_2[7]
port 447 nsew signal output
rlabel metal3 s 0 117678 2226 117738 6 y_r_2[8]
port 448 nsew signal output
rlabel metal2 s 67652 0 67680 2252 6 y_r_2[9]
port 449 nsew signal output
rlabel metal2 s 12912 0 12940 2796 6 y_r_3[0]
port 450 nsew signal output
rlabel metal2 s 25148 116884 25176 120000 6 y_r_3[10]
port 451 nsew signal output
rlabel metal3 s 118110 78918 120000 78978 6 y_r_3[11]
port 452 nsew signal output
rlabel metal2 s 112088 117422 112116 120000 6 y_r_3[12]
port 453 nsew signal output
rlabel metal2 s 48332 0 48360 2252 6 y_r_3[13]
port 454 nsew signal output
rlabel metal3 s 0 29278 386 29338 6 y_r_3[14]
port 455 nsew signal output
rlabel metal3 s 0 718 2226 778 6 y_r_3[15]
port 456 nsew signal output
rlabel metal2 s 95988 0 96016 2252 6 y_r_3[16]
port 457 nsew signal output
rlabel metal2 s 79888 117156 79916 120000 6 y_r_3[1]
port 458 nsew signal output
rlabel metal2 s 92124 0 92152 2796 6 y_r_3[2]
port 459 nsew signal output
rlabel metal2 s 38672 0 38700 2252 6 y_r_3[3]
port 460 nsew signal output
rlabel metal2 s 5828 0 5856 2796 6 y_r_3[4]
port 461 nsew signal output
rlabel metal3 s 117374 2758 120000 2818 6 y_r_3[5]
port 462 nsew signal output
rlabel metal3 s 118110 37438 120000 37498 6 y_r_3[6]
port 463 nsew signal output
rlabel metal2 s 25792 117156 25820 120000 6 y_r_3[7]
port 464 nsew signal output
rlabel metal3 s 117834 114278 120000 114338 6 y_r_3[8]
port 465 nsew signal output
rlabel metal3 s 0 13638 754 13698 6 y_r_3[9]
port 466 nsew signal output
rlabel metal3 s 0 87078 1490 87138 6 y_r_4[0]
port 467 nsew signal output
rlabel metal3 s 0 83678 386 83738 6 y_r_4[10]
port 468 nsew signal output
rlabel metal2 s 5184 0 5212 2252 6 y_r_4[11]
port 469 nsew signal output
rlabel metal3 s 0 11598 754 11658 6 y_r_4[12]
port 470 nsew signal output
rlabel metal3 s 117834 68718 120000 68778 6 y_r_4[13]
port 471 nsew signal output
rlabel metal2 s 70228 0 70256 1170 6 y_r_4[14]
port 472 nsew signal output
rlabel metal2 s 72804 117156 72832 120000 6 y_r_4[15]
port 473 nsew signal output
rlabel metal2 s 102428 117156 102456 120000 6 y_r_4[16]
port 474 nsew signal output
rlabel metal3 s 0 116998 2778 117058 6 y_r_4[1]
port 475 nsew signal output
rlabel metal3 s 0 40838 1490 40898 6 y_r_4[2]
port 476 nsew signal output
rlabel metal3 s 117834 78238 120000 78298 6 y_r_4[3]
port 477 nsew signal output
rlabel metal2 s 106936 117428 106964 120000 6 y_r_4[4]
port 478 nsew signal output
rlabel metal3 s 0 58518 754 58578 6 y_r_4[5]
port 479 nsew signal output
rlabel metal3 s 118110 100678 120000 100738 6 y_r_4[6]
port 480 nsew signal output
rlabel metal3 s 118110 42878 120000 42938 6 y_r_4[7]
port 481 nsew signal output
rlabel metal2 s 83752 0 83780 2252 6 y_r_4[8]
port 482 nsew signal output
rlabel metal2 s 92768 117156 92796 120000 6 y_r_4[9]
port 483 nsew signal output
rlabel metal2 s 21284 117156 21312 120000 6 y_r_5[0]
port 484 nsew signal output
rlabel metal2 s 37384 0 37412 2252 6 y_r_5[10]
port 485 nsew signal output
rlabel metal3 s 118110 77558 120000 77618 6 y_r_5[11]
port 486 nsew signal output
rlabel metal2 s 98564 0 98592 960 6 y_r_5[12]
port 487 nsew signal output
rlabel metal3 s 117834 38118 120000 38178 6 y_r_5[13]
port 488 nsew signal output
rlabel metal3 s 0 53758 1490 53818 6 y_r_5[14]
port 489 nsew signal output
rlabel metal3 s 118110 4798 120000 4858 6 y_r_5[15]
port 490 nsew signal output
rlabel metal2 s 19352 0 19380 2796 6 y_r_5[16]
port 491 nsew signal output
rlabel metal2 s 59924 0 59952 2796 6 y_r_5[1]
port 492 nsew signal output
rlabel metal3 s 118110 55118 120000 55178 6 y_r_5[2]
port 493 nsew signal output
rlabel metal2 s 89548 117428 89576 120000 6 y_r_5[3]
port 494 nsew signal output
rlabel metal3 s 117834 112918 120000 112978 6 y_r_5[4]
port 495 nsew signal output
rlabel metal3 s 117834 5478 120000 5538 6 y_r_5[5]
port 496 nsew signal output
rlabel metal2 s 9692 0 9720 2252 6 y_r_5[6]
port 497 nsew signal output
rlabel metal3 s 118110 71438 120000 71498 6 y_r_5[7]
port 498 nsew signal output
rlabel metal2 s 2608 0 2636 1170 6 y_r_5[8]
port 499 nsew signal output
rlabel metal3 s 118110 115638 120000 115698 6 y_r_5[9]
port 500 nsew signal output
rlabel metal2 s 85684 117156 85712 120000 6 y_r_6[0]
port 501 nsew signal output
rlabel metal3 s 117834 14318 120000 14378 6 y_r_6[10]
port 502 nsew signal output
rlabel metal2 s 82464 117156 82492 120000 6 y_r_6[11]
port 503 nsew signal output
rlabel metal2 s 80532 0 80560 552 6 y_r_6[12]
port 504 nsew signal output
rlabel metal3 s 0 30638 846 30698 6 y_r_6[13]
port 505 nsew signal output
rlabel metal2 s 79888 0 79916 1170 6 y_r_6[14]
port 506 nsew signal output
rlabel metal2 s 32 0 60 1232 6 y_r_6[15]
port 507 nsew signal output
rlabel metal2 s 94056 0 94084 2252 6 y_r_6[16]
port 508 nsew signal output
rlabel metal3 s 0 52398 846 52458 6 y_r_6[1]
port 509 nsew signal output
rlabel metal3 s 0 1398 1122 1458 6 y_r_6[2]
port 510 nsew signal output
rlabel metal2 s 30944 117156 30972 120000 6 y_r_6[3]
port 511 nsew signal output
rlabel metal3 s 0 34718 386 34778 6 y_r_6[4]
port 512 nsew signal output
rlabel metal2 s 24504 0 24532 2252 6 y_r_6[5]
port 513 nsew signal output
rlabel metal2 s 8404 0 8432 2252 6 y_r_6[6]
port 514 nsew signal output
rlabel metal2 s 61212 117156 61240 120000 6 y_r_6[7]
port 515 nsew signal output
rlabel metal2 s 34808 117156 34836 120000 6 y_r_6[8]
port 516 nsew signal output
rlabel metal2 s 63788 0 63816 2252 6 y_r_6[9]
port 517 nsew signal output
rlabel metal2 s 81176 119870 81204 120000 6 y_r_7[0]
port 518 nsew signal output
rlabel metal3 s 117834 32678 120000 32738 6 y_r_7[10]
port 519 nsew signal output
rlabel metal3 s 0 77558 662 77618 6 y_r_7[11]
port 520 nsew signal output
rlabel metal3 s 117098 93878 120000 93938 6 y_r_7[12]
port 521 nsew signal output
rlabel metal2 s 26436 0 26464 2796 6 y_r_7[13]
port 522 nsew signal output
rlabel metal2 s 45756 0 45784 2252 6 y_r_7[14]
port 523 nsew signal output
rlabel metal3 s 0 8198 1490 8258 6 y_r_7[15]
port 524 nsew signal output
rlabel metal3 s 117374 89118 120000 89178 6 y_r_7[16]
port 525 nsew signal output
rlabel metal2 s 70872 0 70900 2252 6 y_r_7[1]
port 526 nsew signal output
rlabel metal2 s 78600 117428 78628 120000 6 y_r_7[2]
port 527 nsew signal output
rlabel metal2 s 77956 117156 77984 120000 6 y_r_7[3]
port 528 nsew signal output
rlabel metal3 s 0 112918 570 112978 6 y_r_7[4]
port 529 nsew signal output
rlabel metal2 s 14200 117156 14228 120000 6 y_r_7[5]
port 530 nsew signal output
rlabel metal2 s 85040 0 85068 688 6 y_r_7[6]
port 531 nsew signal output
rlabel metal3 s 0 26558 386 26618 6 y_r_7[7]
port 532 nsew signal output
rlabel metal3 s 0 102038 662 102098 6 y_r_7[8]
port 533 nsew signal output
rlabel metal3 s 117834 57838 120000 57898 6 y_r_7[9]
port 534 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 26635846
string GDS_FILE /home/icpedia/Desktop/OpenLane/designs/fft_dit/runs/assignment/RUN_2025.08.22_00.24.08/results/signoff/fft_dit.magic.gds
string GDS_START 940018
<< end >>

