* NGSPICE file created from fft_dit.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt fft_dit clk enable finish rst vccd1 vssd1 x_i_0[0] x_i_0[10] x_i_0[11] x_i_0[12]
+ x_i_0[13] x_i_0[14] x_i_0[15] x_i_0[1] x_i_0[2] x_i_0[3] x_i_0[4] x_i_0[5] x_i_0[6]
+ x_i_0[7] x_i_0[8] x_i_0[9] x_i_1[0] x_i_1[10] x_i_1[11] x_i_1[12] x_i_1[13] x_i_1[14]
+ x_i_1[15] x_i_1[1] x_i_1[2] x_i_1[3] x_i_1[4] x_i_1[5] x_i_1[6] x_i_1[7] x_i_1[8]
+ x_i_1[9] x_i_2[0] x_i_2[10] x_i_2[11] x_i_2[12] x_i_2[13] x_i_2[14] x_i_2[15] x_i_2[1]
+ x_i_2[2] x_i_2[3] x_i_2[4] x_i_2[5] x_i_2[6] x_i_2[7] x_i_2[8] x_i_2[9] x_i_3[0]
+ x_i_3[10] x_i_3[11] x_i_3[12] x_i_3[13] x_i_3[14] x_i_3[15] x_i_3[1] x_i_3[2] x_i_3[3]
+ x_i_3[4] x_i_3[5] x_i_3[6] x_i_3[7] x_i_3[8] x_i_3[9] x_i_4[0] x_i_4[10] x_i_4[11]
+ x_i_4[12] x_i_4[13] x_i_4[14] x_i_4[15] x_i_4[1] x_i_4[2] x_i_4[3] x_i_4[4] x_i_4[5]
+ x_i_4[6] x_i_4[7] x_i_4[8] x_i_4[9] x_i_5[0] x_i_5[10] x_i_5[11] x_i_5[12] x_i_5[13]
+ x_i_5[14] x_i_5[15] x_i_5[1] x_i_5[2] x_i_5[3] x_i_5[4] x_i_5[5] x_i_5[6] x_i_5[7]
+ x_i_5[8] x_i_5[9] x_i_6[0] x_i_6[10] x_i_6[11] x_i_6[12] x_i_6[13] x_i_6[14] x_i_6[15]
+ x_i_6[1] x_i_6[2] x_i_6[3] x_i_6[4] x_i_6[5] x_i_6[6] x_i_6[7] x_i_6[8] x_i_6[9]
+ x_i_7[0] x_i_7[10] x_i_7[11] x_i_7[12] x_i_7[13] x_i_7[14] x_i_7[15] x_i_7[1] x_i_7[2]
+ x_i_7[3] x_i_7[4] x_i_7[5] x_i_7[6] x_i_7[7] x_i_7[8] x_i_7[9] x_r_0[0] x_r_0[10]
+ x_r_0[11] x_r_0[12] x_r_0[13] x_r_0[14] x_r_0[15] x_r_0[1] x_r_0[2] x_r_0[3] x_r_0[4]
+ x_r_0[5] x_r_0[6] x_r_0[7] x_r_0[8] x_r_0[9] x_r_1[0] x_r_1[10] x_r_1[11] x_r_1[12]
+ x_r_1[13] x_r_1[14] x_r_1[15] x_r_1[1] x_r_1[2] x_r_1[3] x_r_1[4] x_r_1[5] x_r_1[6]
+ x_r_1[7] x_r_1[8] x_r_1[9] x_r_2[0] x_r_2[10] x_r_2[11] x_r_2[12] x_r_2[13] x_r_2[14]
+ x_r_2[15] x_r_2[1] x_r_2[2] x_r_2[3] x_r_2[4] x_r_2[5] x_r_2[6] x_r_2[7] x_r_2[8]
+ x_r_2[9] x_r_3[0] x_r_3[10] x_r_3[11] x_r_3[12] x_r_3[13] x_r_3[14] x_r_3[15] x_r_3[1]
+ x_r_3[2] x_r_3[3] x_r_3[4] x_r_3[5] x_r_3[6] x_r_3[7] x_r_3[8] x_r_3[9] x_r_4[0]
+ x_r_4[10] x_r_4[11] x_r_4[12] x_r_4[13] x_r_4[14] x_r_4[15] x_r_4[1] x_r_4[2] x_r_4[3]
+ x_r_4[4] x_r_4[5] x_r_4[6] x_r_4[7] x_r_4[8] x_r_4[9] x_r_5[0] x_r_5[10] x_r_5[11]
+ x_r_5[12] x_r_5[13] x_r_5[14] x_r_5[15] x_r_5[1] x_r_5[2] x_r_5[3] x_r_5[4] x_r_5[5]
+ x_r_5[6] x_r_5[7] x_r_5[8] x_r_5[9] x_r_6[0] x_r_6[10] x_r_6[11] x_r_6[12] x_r_6[13]
+ x_r_6[14] x_r_6[15] x_r_6[1] x_r_6[2] x_r_6[3] x_r_6[4] x_r_6[5] x_r_6[6] x_r_6[7]
+ x_r_6[8] x_r_6[9] x_r_7[0] x_r_7[10] x_r_7[11] x_r_7[12] x_r_7[13] x_r_7[14] x_r_7[15]
+ x_r_7[1] x_r_7[2] x_r_7[3] x_r_7[4] x_r_7[5] x_r_7[6] x_r_7[7] x_r_7[8] x_r_7[9]
+ y_i_0[0] y_i_0[10] y_i_0[11] y_i_0[12] y_i_0[13] y_i_0[14] y_i_0[15] y_i_0[16] y_i_0[1]
+ y_i_0[2] y_i_0[3] y_i_0[4] y_i_0[5] y_i_0[6] y_i_0[7] y_i_0[8] y_i_0[9] y_i_1[0]
+ y_i_1[10] y_i_1[11] y_i_1[12] y_i_1[13] y_i_1[14] y_i_1[15] y_i_1[16] y_i_1[1] y_i_1[2]
+ y_i_1[3] y_i_1[4] y_i_1[5] y_i_1[6] y_i_1[7] y_i_1[8] y_i_1[9] y_i_2[0] y_i_2[10]
+ y_i_2[11] y_i_2[12] y_i_2[13] y_i_2[14] y_i_2[15] y_i_2[16] y_i_2[1] y_i_2[2] y_i_2[3]
+ y_i_2[4] y_i_2[5] y_i_2[6] y_i_2[7] y_i_2[8] y_i_2[9] y_i_3[0] y_i_3[10] y_i_3[11]
+ y_i_3[12] y_i_3[13] y_i_3[14] y_i_3[15] y_i_3[16] y_i_3[1] y_i_3[2] y_i_3[3] y_i_3[4]
+ y_i_3[5] y_i_3[6] y_i_3[7] y_i_3[8] y_i_3[9] y_i_4[0] y_i_4[10] y_i_4[11] y_i_4[12]
+ y_i_4[13] y_i_4[14] y_i_4[15] y_i_4[16] y_i_4[1] y_i_4[2] y_i_4[3] y_i_4[4] y_i_4[5]
+ y_i_4[6] y_i_4[7] y_i_4[8] y_i_4[9] y_i_5[0] y_i_5[10] y_i_5[11] y_i_5[12] y_i_5[13]
+ y_i_5[14] y_i_5[15] y_i_5[16] y_i_5[1] y_i_5[2] y_i_5[3] y_i_5[4] y_i_5[5] y_i_5[6]
+ y_i_5[7] y_i_5[8] y_i_5[9] y_i_6[0] y_i_6[10] y_i_6[11] y_i_6[12] y_i_6[13] y_i_6[14]
+ y_i_6[15] y_i_6[16] y_i_6[1] y_i_6[2] y_i_6[3] y_i_6[4] y_i_6[5] y_i_6[6] y_i_6[7]
+ y_i_6[8] y_i_6[9] y_i_7[0] y_i_7[10] y_i_7[11] y_i_7[12] y_i_7[13] y_i_7[14] y_i_7[15]
+ y_i_7[16] y_i_7[1] y_i_7[2] y_i_7[3] y_i_7[4] y_i_7[5] y_i_7[6] y_i_7[7] y_i_7[8]
+ y_i_7[9] y_r_0[0] y_r_0[10] y_r_0[11] y_r_0[12] y_r_0[13] y_r_0[14] y_r_0[15] y_r_0[16]
+ y_r_0[1] y_r_0[2] y_r_0[3] y_r_0[4] y_r_0[5] y_r_0[6] y_r_0[7] y_r_0[8] y_r_0[9]
+ y_r_1[0] y_r_1[10] y_r_1[11] y_r_1[12] y_r_1[13] y_r_1[14] y_r_1[15] y_r_1[16] y_r_1[1]
+ y_r_1[2] y_r_1[3] y_r_1[4] y_r_1[5] y_r_1[6] y_r_1[7] y_r_1[8] y_r_1[9] y_r_2[0]
+ y_r_2[10] y_r_2[11] y_r_2[12] y_r_2[13] y_r_2[14] y_r_2[15] y_r_2[16] y_r_2[1] y_r_2[2]
+ y_r_2[3] y_r_2[4] y_r_2[5] y_r_2[6] y_r_2[7] y_r_2[8] y_r_2[9] y_r_3[0] y_r_3[10]
+ y_r_3[11] y_r_3[12] y_r_3[13] y_r_3[14] y_r_3[15] y_r_3[16] y_r_3[1] y_r_3[2] y_r_3[3]
+ y_r_3[4] y_r_3[5] y_r_3[6] y_r_3[7] y_r_3[8] y_r_3[9] y_r_4[0] y_r_4[10] y_r_4[11]
+ y_r_4[12] y_r_4[13] y_r_4[14] y_r_4[15] y_r_4[16] y_r_4[1] y_r_4[2] y_r_4[3] y_r_4[4]
+ y_r_4[5] y_r_4[6] y_r_4[7] y_r_4[8] y_r_4[9] y_r_5[0] y_r_5[10] y_r_5[11] y_r_5[12]
+ y_r_5[13] y_r_5[14] y_r_5[15] y_r_5[16] y_r_5[1] y_r_5[2] y_r_5[3] y_r_5[4] y_r_5[5]
+ y_r_5[6] y_r_5[7] y_r_5[8] y_r_5[9] y_r_6[0] y_r_6[10] y_r_6[11] y_r_6[12] y_r_6[13]
+ y_r_6[14] y_r_6[15] y_r_6[16] y_r_6[1] y_r_6[2] y_r_6[3] y_r_6[4] y_r_6[5] y_r_6[6]
+ y_r_6[7] y_r_6[8] y_r_6[9] y_r_7[0] y_r_7[10] y_r_7[11] y_r_7[12] y_r_7[13] y_r_7[14]
+ y_r_7[15] y_r_7[16] y_r_7[1] y_r_7[2] y_r_7[3] y_r_7[4] y_r_7[5] y_r_7[6] y_r_7[7]
+ y_r_7[8] y_r_7[9]
XFILLER_140_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09671_ _09670_/Y _15553_/Q _09669_/B vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07534__A1 input109/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08622_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08553_ _08549_/B _08553_/B vssd1 vssd1 vccd1 vccd1 _08553_/X sky130_fd_sc_hd__and2b_1
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11094__A1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _15512_/Q input28/X _07536_/S vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08484_ _08484_/A _08499_/C vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__xnor2_1
XFILLER_211_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ _15546_/Q _07435_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07436_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14446__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ _15502_/Q _15486_/Q vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__and2_1
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _15376_/Q _15360_/Q vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__or2b_1
XFILLER_50_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14181__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09275__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13509__B _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07773__A1 _07773_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _09938_/A _09946_/A vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ _15218_/Q _09971_/B vssd1 vssd1 vccd1 vccd1 _09869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ _11901_/A _11901_/B _11901_/C vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__a21o_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input127_A x_i_7[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12880_ _12730_/A _12835_/Y _12837_/B vssd1 vssd1 vccd1 vccd1 _13018_/B sky130_fd_sc_hd__o21ai_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11831_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _12415_/B sky130_fd_sc_hd__nand2_2
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14550_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14550_/Y sky130_fd_sc_hd__inv_2
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11808_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__nor2_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13501_ _13501_/A vssd1 vssd1 vccd1 vccd1 _15640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10713_ _10713_/A _11014_/A vssd1 vssd1 vccd1 vccd1 _15051_/D sky130_fd_sc_hd__xor2_4
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__buf_6
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _12144_/A _12008_/A _11692_/C vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__a21oi_1
XFILLER_158_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14356__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07669__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ _13432_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__or2_1
XANTENNA_input92_A x_i_5[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10644_ _10972_/A _10644_/B vssd1 vssd1 vccd1 vccd1 _15039_/D sky130_fd_sc_hd__xnor2_4
XFILLER_42_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08354__A _15726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _13362_/A _13362_/B _13362_/C vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__a21o_1
X_10575_ _10575_/A vssd1 vssd1 vccd1 vccd1 _15033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ _15346_/CLK _15102_/D _14143_/Y vssd1 vssd1 vccd1 vccd1 _15102_/Q sky130_fd_sc_hd__dfrtp_1
X_12314_ _12511_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__xnor2_4
XFILLER_6_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13294_ _13737_/B _13295_/B _13293_/Y _13217_/Y vssd1 vssd1 vccd1 vccd1 _13294_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1068 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15033_ _15483_/CLK _15033_/D _14070_/Y vssd1 vssd1 vccd1 vccd1 _15033_/Q sky130_fd_sc_hd__dfrtp_1
X_12245_ _12247_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14091__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12176_ _12240_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__and2_1
XFILLER_190_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12323__B _12323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11127_/A _11127_/B _11127_/C vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__nor3_1
XFILLER_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11058_ _14930_/Q _14996_/Q vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output513_A output513/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07516__A1 _07516_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10009_ _10009_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _14937_/D sky130_fd_sc_hd__xnor2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14817_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15797_ _15799_/CLK _15797_/D _14877_/Y vssd1 vssd1 vccd1 vccd1 _15797_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater663_A _14753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14748_ _14750_/A vssd1 vssd1 vccd1 vccd1 _14748_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater830_A input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14266__A _14269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14679_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15800__D _15800_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_475 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07579__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__B _15480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__A1 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput401 _10797_/Y vssd1 vssd1 vccd1 vccd1 y_r_0[14] sky130_fd_sc_hd__buf_2
Xoutput412 output412/A vssd1 vssd1 vccd1 vccd1 y_r_0[9] sky130_fd_sc_hd__buf_2
Xoutput423 _15580_/Q vssd1 vssd1 vccd1 vccd1 y_r_1[3] sky130_fd_sc_hd__buf_2
XFILLER_160_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput434 output434/A vssd1 vssd1 vccd1 vccd1 y_r_2[13] sky130_fd_sc_hd__buf_2
XANTENNA__09807__B _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput445 output445/A vssd1 vssd1 vccd1 vccd1 y_r_2[8] sky130_fd_sc_hd__buf_2
Xoutput456 _15596_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[2] sky130_fd_sc_hd__buf_2
Xoutput467 output467/A vssd1 vssd1 vccd1 vccd1 y_r_4[12] sky130_fd_sc_hd__buf_2
Xoutput478 _11272_/X vssd1 vssd1 vccd1 vccd1 y_r_4[7] sky130_fd_sc_hd__buf_2
XFILLER_114_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput489 _15611_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[1] sky130_fd_sc_hd__buf_2
XANTENNA__07755__A1 _07755_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ _11584_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08074_/C sky130_fd_sc_hd__xor2_1
XFILLER_80_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09723_ _09840_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _15717_/D sky130_fd_sc_hd__xnor2_1
XFILLER_45_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09654_ _09654_/A _09654_/B _09654_/C vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__or3_1
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10688__B _15279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _12654_/A _08500_/Y _08570_/B _12627_/A _08604_/X vssd1 vssd1 vccd1 vccd1
+ _08605_/X sky130_fd_sc_hd__o221a_1
X_09585_ _09793_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _09590_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08158__B _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _13030_/C _08550_/A _08536_/C vssd1 vssd1 vccd1 vccd1 _08546_/B sky130_fd_sc_hd__or3_2
XFILLER_208_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08467_ _08587_/A _08587_/B _08466_/X vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__a21oi_2
XFILLER_169_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14176__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13080__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__A0 _15420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07418_ _15554_/Q input55/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07419_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ _15045_/Q vssd1 vssd1 vccd1 vccd1 _13201_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_93_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ _10360_/A _10360_/B _10480_/A vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__and3_1
XFILLER_163_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _15374_/Q _15358_/Q vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__nor2_1
XFILLER_163_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10291_ _10291_/A _11430_/A vssd1 vssd1 vccd1 vccd1 _15774_/D sky130_fd_sc_hd__xnor2_1
X_12030_ _12030_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__or2_1
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__A1 _07746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input244_A x_r_7[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_862 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13981_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13981_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15720_ _15722_/CLK _15720_/D _14796_/Y vssd1 vssd1 vccd1 vccd1 _15720_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _13203_/A _12933_/B _13006_/A _12931_/X vssd1 vssd1 vccd1 vccd1 _12934_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15689_/CLK _15651_/D _14724_/Y vssd1 vssd1 vccd1 vccd1 _15651_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ _12863_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12951_/C sky130_fd_sc_hd__xor2_1
XFILLER_61_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14602_/Y sky130_fd_sc_hd__inv_2
X_11814_ _11814_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11815_/B sky130_fd_sc_hd__or2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15680_/CLK _15582_/D _14651_/Y vssd1 vssd1 vccd1 vccd1 _15582_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12794_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__xnor2_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14533_/Y sky130_fd_sc_hd__inv_2
X_11745_ _11833_/A _11833_/B vssd1 vssd1 vccd1 vccd1 _11834_/A sky130_fd_sc_hd__xnor2_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14086__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14464_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14464_/Y sky130_fd_sc_hd__inv_2
X_11676_ _11676_/A _11775_/A vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__xnor2_1
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12318__B _12323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _13416_/A _15052_/Q vssd1 vssd1 vccd1 vccd1 _13417_/A sky130_fd_sc_hd__and2_1
XFILLER_186_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10627_ _10585_/B _10625_/B _10626_/Y vssd1 vssd1 vccd1 vccd1 _10628_/B sky130_fd_sc_hd__o21ai_1
XFILLER_128_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14395_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14814__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13346_ _15768_/Q _13572_/A vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__xor2_1
XFILLER_143_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10558_ _10558_/A _10558_/B _10612_/A vssd1 vssd1 vccd1 vccd1 _10558_/X sky130_fd_sc_hd__and3_1
XFILLER_182_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output463_A output463/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13277_ _13205_/A _13277_/B vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__and2b_1
X_10489_ _10496_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__nand2_1
X_15016_ _15435_/CLK _15016_/D _14052_/Y vssd1 vssd1 vccd1 vccd1 _15016_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__inv_2
XFILLER_155_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13149__B _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ _15737_/Q vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__inv_2
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater904 input215/X vssd1 vssd1 vccd1 vccd1 _07712_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07862__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater915 input198/X vssd1 vssd1 vccd1 vccd1 _07844_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater926 repeater927/X vssd1 vssd1 vccd1 vccd1 _07706_/A1 sky130_fd_sc_hd__buf_4
XFILLER_110_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater780_A repeater781/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater937 input164/X vssd1 vssd1 vccd1 vccd1 _07816_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater948 input150/X vssd1 vssd1 vccd1 vccd1 _07746_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater959 input136/X vssd1 vssd1 vccd1 vccd1 _07872_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09370_ _09368_/A _09368_/B _09369_/X vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__a21o_1
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08321_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ _11832_/A _08292_/B _08288_/A _08252_/D vssd1 vssd1 vccd1 vccd1 _08288_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_166_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08183_ _15015_/Q vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__buf_6
XFILLER_158_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _14904_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_20_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14724__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12244__A _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput264 _11088_/X vssd1 vssd1 vccd1 vccd1 y_i_0[13] sky130_fd_sc_hd__buf_2
XFILLER_173_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07728__A1 input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput275 output275/A vssd1 vssd1 vccd1 vccd1 y_i_0[8] sky130_fd_sc_hd__buf_2
XFILLER_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput286 _15645_/Q vssd1 vssd1 vccd1 vccd1 y_i_1[2] sky130_fd_sc_hd__buf_2
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput297 _10941_/X vssd1 vssd1 vccd1 vccd1 y_i_2[12] sky130_fd_sc_hd__buf_2
XFILLER_181_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07967_ _15775_/Q vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__inv_2
XFILLER_210_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _09706_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__nand2_2
XFILLER_210_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09272__B _15492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07898_ _15318_/Q input138/X _07900_/S vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _15564_/Q _15544_/Q vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__and2b_1
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07900__A1 input131/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _15436_/Q _15420_/Q vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__xnor2_2
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08519_ _12688_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08525_/A sky130_fd_sc_hd__nor2_1
XFILLER_180_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09499_ _15527_/Q _15511_/Q _09498_/B vssd1 vssd1 vccd1 vccd1 _09499_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11530_ _11530_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__xnor2_1
XFILLER_168_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11461_ _11509_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11462_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input194_A x_r_3[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14634__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200_ _13201_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _13274_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ _10412_/A _10412_/B _10412_/C vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__or3_1
XFILLER_171_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14180_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14180_/Y sky130_fd_sc_hd__inv_2
X_11392_ _11392_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _15727_/D sky130_fd_sc_hd__xnor2_1
XFILLER_164_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13131_/A _13131_/B vssd1 vssd1 vccd1 vccd1 _13703_/B sky130_fd_sc_hd__nor2_4
X_10343_ _15129_/Q _15162_/Q vssd1 vssd1 vccd1 vccd1 _10343_/X sky130_fd_sc_hd__and2_1
XFILLER_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input55_A x_i_3[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _13702_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__nor2_1
X_10274_ _10274_/A _10274_/B _11421_/A vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__and3_1
XFILLER_2_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _11935_/A _11935_/B _11933_/A _11932_/A vssd1 vssd1 vccd1 vccd1 _12014_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_2_0_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15615__D _15615_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13964_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13964_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15703_ _15770_/CLK _15703_/D _14778_/Y vssd1 vssd1 vccd1 vccd1 _15703_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12915_ _12841_/A _13669_/B _12914_/Y vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__a21boi_4
XFILLER_59_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13895_ _13895_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _15062_/D sky130_fd_sc_hd__xnor2_1
XFILLER_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14809__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output309_A output309/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15634_ _15784_/CLK _15634_/D _14706_/Y vssd1 vssd1 vccd1 vccd1 _15634_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ _13537_/A _12846_/B vssd1 vssd1 vccd1 vccd1 _15629_/D sky130_fd_sc_hd__xnor2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _15592_/CLK _15565_/D _14632_/Y vssd1 vssd1 vccd1 vccd1 _15565_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12777_ _12777_/A _12777_/B _12777_/C vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__and3_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A _11233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07655__A0 _15438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14516_/Y sky130_fd_sc_hd__inv_2
X_11728_ _11728_/A _12390_/A vssd1 vssd1 vccd1 vccd1 _11728_/Y sky130_fd_sc_hd__xnor2_1
X_15496_ _15569_/CLK _15496_/D _14559_/Y vssd1 vssd1 vccd1 vccd1 _15496_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14447_/Y sky130_fd_sc_hd__inv_2
X_11659_ _11606_/B _11659_/B vssd1 vssd1 vccd1 vccd1 _11659_/X sky130_fd_sc_hd__and2b_1
XFILLER_175_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_940 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14544__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08604__C1 _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14378_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10791__B _15788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329_ _13374_/A _13329_/B vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__xnor2_1
XFILLER_143_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_142_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08870_ _08945_/A _08867_/B _08869_/X vssd1 vssd1 vccd1 vccd1 _08871_/B sky130_fd_sc_hd__a21o_1
Xrepeater701 _07695_/S vssd1 vssd1 vccd1 vccd1 _07697_/S sky130_fd_sc_hd__buf_6
X_07821_ _07821_/A vssd1 vssd1 vccd1 vccd1 _15357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater712 _15708_/Q vssd1 vssd1 vccd1 vccd1 output386/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater723 _15692_/Q vssd1 vssd1 vccd1 vccd1 output352/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater734 _15672_/Q vssd1 vssd1 vccd1 vccd1 output314/A sky130_fd_sc_hd__clkbuf_2
Xrepeater745 repeater746/X vssd1 vssd1 vccd1 vccd1 output280/A sky130_fd_sc_hd__buf_4
X_07752_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07795_/S sky130_fd_sc_hd__buf_6
Xrepeater756 _15646_/Q vssd1 vssd1 vccd1 vccd1 repeater756/X sky130_fd_sc_hd__buf_4
Xrepeater767 _15631_/Q vssd1 vssd1 vccd1 vccd1 output527/A sky130_fd_sc_hd__clkbuf_2
Xrepeater778 repeater779/X vssd1 vssd1 vccd1 vccd1 output496/A sky130_fd_sc_hd__buf_6
XFILLER_37_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater789 _15603_/Q vssd1 vssd1 vccd1 vccd1 output463/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07683_ _15424_/Q input181/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_898 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14719__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13623__A _15377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _15529_/Q _15513_/Q vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__nand2_1
XFILLER_164_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ _09353_/A vssd1 vssd1 vccd1 vccd1 _15136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08304_ _08304_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__and2_1
X_09284_ _09284_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _15121_/D sky130_fd_sc_hd__xnor2_1
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__xor2_2
XFILLER_119_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14454__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_798 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07767__S _07795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08166_ _11906_/A _11707_/A vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10973__B_N _15270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08452__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08097_ _11898_/A _08097_/B vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__xnor2_2
XFILLER_162_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08374__A1 _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ _15370_/Q _15354_/Q vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__xnor2_2
XFILLER_47_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10222__A _15075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_887 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ _14970_/Q _14904_/Q vssd1 vssd1 vccd1 vccd1 _11143_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14629__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12700_ _12700_/A _13529_/B vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__or2_1
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13680_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__inv_2
X_10892_ _14960_/Q _14894_/Q vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input207_A x_r_4[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__A_N _15466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13252__B _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _12630_/A _12810_/A _08654_/B _12921_/A _13012_/A vssd1 vssd1 vccd1 vccd1
+ _12635_/A sky130_fd_sc_hd__o2111a_1
XFILLER_34_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _15460_/CLK _15350_/D _14405_/Y vssd1 vssd1 vccd1 vccd1 _15350_/Q sky130_fd_sc_hd__dfrtp_1
X_12562_ _15737_/Q _12219_/B _12561_/X vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14301_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14301_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11513_ _11678_/A _11658_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__and3b_1
XFILLER_184_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15281_ _15400_/CLK _15281_/D _14332_/Y vssd1 vssd1 vccd1 vccd1 _15281_/Q sky130_fd_sc_hd__dfrtp_2
X_12493_ _12493_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__xor2_1
XANTENNA__14364__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07677__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__inv_2
X_11444_ _11527_/A _11527_/B vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__xor2_1
XFILLER_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14163_/Y sky130_fd_sc_hd__inv_2
X_11375_ _11375_/A _11375_/B _11375_/C vssd1 vssd1 vccd1 vccd1 _11377_/A sky130_fd_sc_hd__nor3_1
XFILLER_3_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13114_ _13147_/A _13146_/A vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10326_ _10459_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _15782_/D sky130_fd_sc_hd__xnor2_4
XFILLER_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__inv_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output259_A output259/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13046_/A _13046_/B vssd1 vssd1 vccd1 vccd1 _13124_/B sky130_fd_sc_hd__nand2_1
X_10257_ _15080_/Q _15245_/Q vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__or2b_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10188_ _15235_/Q _15070_/Q vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__or2b_1
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output426_A output426/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11228__A _15033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14996_ _15498_/CLK _14996_/D _14030_/Y vssd1 vssd1 vccd1 vccd1 _14996_/Q sky130_fd_sc_hd__dfrtp_1
X_13947_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13947_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14539__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater576_A repeater577/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13878_ _15335_/Q _15319_/Q _13877_/B vssd1 vssd1 vccd1 vccd1 _13878_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15617_ _15617_/CLK _15617_/D _14688_/Y vssd1 vssd1 vccd1 vccd1 _15617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ _12882_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07628__A0 _15451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15548_ _15563_/CLK _15548_/D _14614_/Y vssd1 vssd1 vccd1 vccd1 _15548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11898__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater910_A input203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15479_ _15542_/CLK _15479_/D _14542_/Y vssd1 vssd1 vccd1 vccd1 _15479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14274__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _08020_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11438_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07587__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _09971_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _14922_/D sky130_fd_sc_hd__xnor2_1
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08922_ _08921_/A _08921_/B _08970_/A vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ _08855_/B _08853_/B vssd1 vssd1 vccd1 vccd1 _15202_/D sky130_fd_sc_hd__nor2_1
XFILLER_112_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07804_ _07804_/A vssd1 vssd1 vccd1 vccd1 _15365_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater542 _10958_/Y vssd1 vssd1 vccd1 vccd1 output300/A sky130_fd_sc_hd__clkbuf_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _15339_/Q _15323_/Q vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__nand2_1
Xrepeater553 _11385_/X vssd1 vssd1 vccd1 vccd1 output435/A sky130_fd_sc_hd__clkbuf_2
Xrepeater564 repeater565/X vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__buf_4
XFILLER_66_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater575 _11332_/X vssd1 vssd1 vccd1 vccd1 output344/A sky130_fd_sc_hd__clkbuf_2
Xrepeater586 repeater587/X vssd1 vssd1 vccd1 vccd1 output261/A sky130_fd_sc_hd__buf_4
X_07735_ _07735_/A vssd1 vssd1 vccd1 vccd1 _15399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater597 _11119_/Y vssd1 vssd1 vccd1 vccd1 output377/A sky130_fd_sc_hd__buf_4
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14449__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07666_ _07666_/A vssd1 vssd1 vccd1 vccd1 _15433_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08447__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10696__B _15280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ _09403_/A _09403_/B _09404_/X vssd1 vssd1 vccd1 vccd1 _15151_/D sky130_fd_sc_hd__a21o_1
XFILLER_77_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07597_ _07597_/A vssd1 vssd1 vccd1 vccd1 _15467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_205_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08166__B _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09336_ _09336_/A _09397_/A vssd1 vssd1 vccd1 vccd1 _15132_/D sky130_fd_sc_hd__xor2_4
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _09266_/A _09266_/C _09266_/B vssd1 vssd1 vccd1 vccd1 _09268_/B sky130_fd_sc_hd__a21oi_1
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14184__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08292_/B _08218_/B vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09198_ _09196_/A _09663_/B _09197_/X vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__a21o_1
XFILLER_135_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08149_ _11906_/A _11707_/A vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__xor2_2
XFILLER_135_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _15744_/Q _11159_/Y _11155_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10111_ _15138_/Q _15303_/Q vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__nand2_1
X_11091_ _15001_/Q _14935_/Q vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input157_A x_r_1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _15208_/Q _15109_/Q vssd1 vssd1 vccd1 vccd1 _10043_/B sky130_fd_sc_hd__nand2_1
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14850_/Y sky130_fd_sc_hd__inv_2
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _13794_/A _13801_/B vssd1 vssd1 vccd1 vccd1 _13801_/X sky130_fd_sc_hd__and2b_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input18_A x_i_0[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ _14781_/A vssd1 vssd1 vccd1 vccd1 _14781_/Y sky130_fd_sc_hd__inv_2
X_11993_ _12144_/A _11692_/C _11992_/Y vssd1 vssd1 vccd1 vccd1 _11994_/C sky130_fd_sc_hd__a21oi_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14359__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A0 _15338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13732_ _14978_/Q _13836_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13732_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10944_ _10944_/A _10950_/A vssd1 vssd1 vccd1 vccd1 _11134_/A sky130_fd_sc_hd__nand2_4
XANTENNA__08357__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13663_ _13663_/A _13663_/B vssd1 vssd1 vccd1 vccd1 _13664_/B sky130_fd_sc_hd__nand2_2
X_10875_ _11109_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__xor2_1
XFILLER_108_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15402_ _15588_/CLK _15402_/D _14460_/Y vssd1 vssd1 vccd1 vccd1 _15402_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12614_/A _12614_/B vssd1 vssd1 vccd1 vccd1 _15690_/D sky130_fd_sc_hd__xnor2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _13594_/A _13594_/B vssd1 vssd1 vccd1 vccd1 _15088_/D sky130_fd_sc_hd__xnor2_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _15782_/CLK _15333_/D _14387_/Y vssd1 vssd1 vccd1 vccd1 _15333_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_200_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _11875_/B _15732_/Q vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__and2b_1
XFILLER_185_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14094__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_132_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15664_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_200_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15264_ _15539_/CLK _15264_/D _14314_/Y vssd1 vssd1 vccd1 vccd1 _15264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12476_ _12460_/A _12602_/B _12604_/A _12475_/Y vssd1 vssd1 vccd1 vccd1 _12488_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output376_A _11117_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14215_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11427_ _11427_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__xnor2_2
X_15195_ _15472_/CLK _15195_/D _14242_/Y vssd1 vssd1 vccd1 vccd1 _15195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _11158_/A _11357_/B _11158_/B vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__a21boi_2
XFILLER_112_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ _10307_/Y _10309_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__and2b_2
XFILLER_141_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13438__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14077_/Y sky130_fd_sc_hd__inv_2
X_11289_ _11289_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11289_/Y sky130_fd_sc_hd__nor2_2
XFILLER_117_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13028_ _13438_/A _13381_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater693_A _08118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07870__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater958_A input137/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14269__A _14269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ _15773_/CLK _14979_/D _14012_/Y vssd1 vssd1 vccd1 vccd1 _14979_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15803__D _15803_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07520_ _15504_/Q input101/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07521_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07451_ _15538_/Q _07451_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07452_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07382_ _15576_/Q input121/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07383_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09121_ _09121_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _15229_/D sky130_fd_sc_hd__xor2_1
XFILLER_202_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15202_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09052_ _09052_/A _09052_/B _13625_/A vssd1 vssd1 vccd1 vccd1 _09054_/A sky130_fd_sc_hd__and3_1
XFILLER_198_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08003_ _08004_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__nor2_1
XFILLER_190_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14732__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09954_ _09953_/A _09953_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__a21o_1
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ _15472_/Q _15456_/Q vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__or2b_1
XFILLER_131_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09885_ _15189_/Q _15222_/Q vssd1 vssd1 vccd1 vccd1 _09885_/Y sky130_fd_sc_hd__nor2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08836_ _08836_/A _08836_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__nor3_1
XFILLER_131_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08767_ _08766_/A _08766_/B _13877_/A vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__o21a_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14179__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _15407_/Q input212/X _07750_/S vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__mux2_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08177__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08698_ _08728_/A _08530_/B _08697_/X vssd1 vssd1 vccd1 vccd1 _12692_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _15441_/Q input246/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07650_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10660_ _15274_/Q _15175_/Q vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__or2_1
XFILLER_15_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ _09319_/A _09386_/A vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__nand2_1
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ _15252_/Q _15285_/Q _10490_/Y _10963_/A vssd1 vssd1 vccd1 vccd1 _10592_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_114_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15761_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12427__A _12439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12244_/A _12328_/Y _12330_/S vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ _12262_/A _12491_/A vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__and2_1
XFILLER_154_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12861__S _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ _14003_/A vssd1 vssd1 vccd1 vccd1 _14000_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11212_ _11212_/A vssd1 vssd1 vccd1 vccd1 _11212_/X sky130_fd_sc_hd__clkbuf_2
X_12192_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__nor2_1
XFILLER_150_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _11143_/A _11143_/B vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__12162__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11074_ _14933_/Q _14999_/Q vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__and2b_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput120 x_i_7[14] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_1
Xinput131 x_r_0[0] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_2
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ _15732_/CLK _14902_/D _13931_/Y vssd1 vssd1 vccd1 vccd1 _14902_/Q sky130_fd_sc_hd__dfrtp_2
Xinput142 x_r_0[5] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__clkbuf_1
X_10025_ _10389_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _14973_/D sky130_fd_sc_hd__xnor2_2
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput153 x_r_1[15] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput164 x_r_2[10] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__clkbuf_1
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 x_r_2[6] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__clkbuf_2
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 x_r_3[1] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_hd__clkbuf_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput197 x_r_4[11] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__clkbuf_2
X_14833_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14833_/Y sky130_fd_sc_hd__inv_2
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14089__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12824__A0 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14764_/Y sky130_fd_sc_hd__inv_2
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08087__A _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _11977_/A _11977_/B vssd1 vssd1 vccd1 vccd1 _12056_/B sky130_fd_sc_hd__nand2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09569__A_N _15435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ _13715_/A _13715_/B vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__nand2_1
X_10927_ _10927_/A vssd1 vssd1 vccd1 vccd1 _10927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14695_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14695_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14817__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13646_ _13669_/A _13646_/B _13646_/C vssd1 vssd1 vccd1 vccd1 _13648_/A sky130_fd_sc_hd__nand3_1
X_10858_ _14955_/Q _15809_/Q vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__or2b_1
XANTENNA_output493_A output493/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_105_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15705_/CLK sky130_fd_sc_hd__clkbuf_16
X_13577_ _15768_/Q _13572_/Y _13575_/X _13576_/X vssd1 vssd1 vccd1 vccd1 _13577_/X
+ sky130_fd_sc_hd__a31o_1
X_10789_ _10787_/X _10795_/A vssd1 vssd1 vccd1 vccd1 _10789_/X sky130_fd_sc_hd__and2b_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater539_A _11243_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15316_ _15575_/CLK _15316_/D _14369_/Y vssd1 vssd1 vccd1 vccd1 _15316_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11241__A _15035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12528_ _12525_/A _12525_/B _12527_/Y vssd1 vssd1 vccd1 vccd1 _12529_/B sky130_fd_sc_hd__a21o_1
XFILLER_145_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15247_ _15764_/CLK _15247_/D _14296_/Y vssd1 vssd1 vccd1 vccd1 _15247_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12459_ _12460_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14552__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater706_A _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ _15663_/CLK _15178_/D _14223_/Y vssd1 vssd1 vccd1 vccd1 _15178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14129_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13168__A _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09670_ _15573_/Q vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _08621_/A _08621_/B vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08552_ _08552_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ _07503_/A vssd1 vssd1 vccd1 vccd1 _15513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11094__A2 _11093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _12871_/A _12780_/A vssd1 vssd1 vccd1 vccd1 _08499_/C sky130_fd_sc_hd__xor2_2
XFILLER_78_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14727__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07485_/S sky130_fd_sc_hd__buf_12
XFILLER_74_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12247__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09104_ _15502_/Q _15486_/Q vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__nor2_1
XFILLER_149_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _15360_/Q _15376_/Q vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__or2b_1
XFILLER_164_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14462__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07775__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09937_ _15229_/Q _15196_/Q vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09868_ _09875_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09971_/B sky130_fd_sc_hd__nand2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _08818_/A _08818_/B _13901_/A vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__a21o_1
XFILLER_133_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A _09799_/B _09799_/C vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nor3_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11829_/B _11829_/C _11829_/A vssd1 vssd1 vccd1 vccd1 _11904_/B sky130_fd_sc_hd__a21o_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11761_ _12178_/A _12055_/A _12038_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12282__B2 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14637__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13500_ _13514_/B _13500_/B vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__and2_1
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10712_/A _10712_/B vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__nor2_4
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14480_/Y sky130_fd_sc_hd__inv_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _12144_/A _12008_/A _11692_/C vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__and3_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13431_ _14920_/Q _13431_/B vssd1 vssd1 vccd1 vccd1 _13432_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08238__B1 _11842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10643_ _10639_/A _10636_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _10644_/B sky130_fd_sc_hd__o21ai_4
XFILLER_167_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input85_A x_i_5[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ _13362_/A _13362_/B _13362_/C vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__and3_1
XFILLER_210_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ _10572_/X _10577_/B vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__and2b_1
XFILLER_194_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15101_ _15375_/CLK _15101_/D _14142_/Y vssd1 vssd1 vccd1 vccd1 _15101_/Q sky130_fd_sc_hd__dfrtp_1
X_12313_ _12329_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12511_/B sky130_fd_sc_hd__xnor2_4
XFILLER_166_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07461__A1 _07461_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ _13217_/A _13722_/B _13292_/Y _13131_/B vssd1 vssd1 vccd1 vccd1 _13293_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__14372__A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07685__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_827 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ _15483_/CLK _15032_/D _14069_/Y vssd1 vssd1 vccd1 vccd1 _15032_/Q sky130_fd_sc_hd__dfrtp_1
X_12244_ _12244_/A vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__inv_2
XFILLER_182_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08370__A _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12175_ _12175_/A _12175_/B _12175_/C vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__nand3_1
XFILLER_3_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11126_ _14964_/Q _14898_/Q vssd1 vssd1 vccd1 vccd1 _11127_/C sky130_fd_sc_hd__and2_1
XFILLER_123_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output339_A _11313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _14930_/Q _14996_/Q vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__or2_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _09966_/B _10006_/B _10007_/Y vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__o21ai_1
XFILLER_209_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output506_A output506/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14816_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14816_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15796_ _15799_/CLK _15796_/D _14876_/Y vssd1 vssd1 vccd1 vccd1 _15796_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11959_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__nand2_1
X_14747_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14747_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12273__B2 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater656_A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14547__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11670__S _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14678_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13629_ _15379_/Q _15363_/Q _13628_/B vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12067__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14282__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput402 _10802_/X vssd1 vssd1 vccd1 vccd1 y_r_0[15] sky130_fd_sc_hd__buf_2
XFILLER_195_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput413 output413/A vssd1 vssd1 vccd1 vccd1 y_r_1[0] sky130_fd_sc_hd__buf_2
Xoutput424 output424/A vssd1 vssd1 vccd1 vccd1 y_r_1[4] sky130_fd_sc_hd__buf_2
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput435 output435/A vssd1 vssd1 vccd1 vccd1 y_r_2[14] sky130_fd_sc_hd__buf_2
XFILLER_126_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput446 _11369_/Y vssd1 vssd1 vccd1 vccd1 y_r_2[9] sky130_fd_sc_hd__buf_2
XFILLER_160_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput457 _15597_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[3] sky130_fd_sc_hd__buf_2
XANTENNA__09095__B _15484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput468 _11294_/X vssd1 vssd1 vccd1 vccd1 y_r_4[13] sky130_fd_sc_hd__buf_2
Xoutput479 output479/A vssd1 vssd1 vccd1 vccd1 y_r_4[8] sky130_fd_sc_hd__buf_2
XFILLER_141_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07983_ _15794_/Q vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__buf_4
XFILLER_86_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _09716_/A _09718_/B _09716_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__a21boi_2
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13626__A _15378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09653_ _15569_/Q _15549_/Q vssd1 vssd1 vccd1 vccd1 _09654_/C sky130_fd_sc_hd__and2b_1
X_08604_ _12627_/A _08570_/B _08530_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08604_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_209_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09584_ _09793_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _15177_/D sky130_fd_sc_hd__xor2_1
XFILLER_83_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ _08728_/A _12688_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08536_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__14457__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08466_ _08466_/A _08466_/B _08466_/C vssd1 vssd1 vccd1 vccd1 _08466_/X sky130_fd_sc_hd__and3_1
XFILLER_51_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07417_ _07417_/A vssd1 vssd1 vccd1 vccd1 _15555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__A1 input192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08397_ _08396_/A _12654_/A _08396_/C vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07443__A1 _07443_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14192__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__B_N _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _13610_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _15110_/D sky130_fd_sc_hd__xor2_1
XFILLER_152_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ _15085_/Q _15250_/Q vssd1 vssd1 vccd1 vccd1 _11430_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13980_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13980_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input237_A x_r_6[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09499__A2 _15511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ _13203_/A _13201_/A _12930_/A _12930_/B vssd1 vssd1 vccd1 vccd1 _12931_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15650_ _15687_/CLK _15650_/D _14723_/Y vssd1 vssd1 vccd1 vccd1 _15650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12862_ _12862_/A _12862_/B vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__xor2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _11814_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__nand2_1
X_14601_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14620_/A sky130_fd_sc_hd__buf_12
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15680_/CLK _15581_/D _14650_/Y vssd1 vssd1 vccd1 vccd1 _15581_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12793_ _12793_/A _12793_/B vssd1 vssd1 vccd1 vccd1 _12794_/B sky130_fd_sc_hd__nor2_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14367__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14532_/Y sky130_fd_sc_hd__inv_2
X_11744_ _11835_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11833_/B sky130_fd_sc_hd__xnor2_1
XFILLER_144_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08365__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14463_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11675_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13414_ _15051_/Q vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__inv_2
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10626_ _15266_/Q _15299_/Q vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__nand2_1
X_14394_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14394_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output289_A _15648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13345_ _13345_/A _13345_/B vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__xnor2_4
XFILLER_154_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10557_ _10557_/A _10565_/A vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__nand2_1
XFILLER_182_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13276_ _13317_/A _13316_/C vssd1 vssd1 vccd1 vccd1 _13280_/A sky130_fd_sc_hd__and2b_1
XFILLER_52_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _15252_/Q _15285_/Q vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__or2b_1
XANTENNA_output456_A _15596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ _15435_/CLK _15015_/D _14051_/Y vssd1 vssd1 vccd1 vccd1 _15015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_1000 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12227_ _12022_/A _12022_/B _12550_/A _12553_/A _12226_/X vssd1 vssd1 vccd1 vccd1
+ _12268_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__14830__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12158_ _12158_/A _12220_/B vssd1 vssd1 vccd1 vccd1 _15587_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11109_ _11109_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_116_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater905 input214/X vssd1 vssd1 vccd1 vccd1 _07714_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_204_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater916 input196/X vssd1 vssd1 vccd1 vccd1 _07848_/A1 sky130_fd_sc_hd__buf_4
XFILLER_96_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12089_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__and3_1
Xrepeater927 input179/X vssd1 vssd1 vccd1 vccd1 repeater927/X sky130_fd_sc_hd__buf_2
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater938 input162/X vssd1 vssd1 vccd1 vccd1 _07753_/A1 sky130_fd_sc_hd__buf_4
Xrepeater949 input149/X vssd1 vssd1 vccd1 vccd1 _07748_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_83_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater773_A _15625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__C_N _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater940_A repeater941/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ _15791_/CLK _15779_/D _14858_/Y vssd1 vssd1 vccd1 vccd1 _15779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14277__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08320_ _12525_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _15577_/D sky130_fd_sc_hd__nand2_1
XFILLER_127_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08251_ _11906_/A _11467_/A vssd1 vssd1 vccd1 vccd1 _08252_/D sky130_fd_sc_hd__or2_1
XFILLER_177_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07673__A1 input243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08182_ _08189_/B _08189_/A vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__and2b_1
XFILLER_119_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14740__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput265 _11095_/Y vssd1 vssd1 vccd1 vccd1 y_i_0[14] sky130_fd_sc_hd__buf_2
XFILLER_160_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput276 output276/A vssd1 vssd1 vccd1 vccd1 y_i_0[9] sky130_fd_sc_hd__buf_2
XFILLER_47_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput287 output287/A vssd1 vssd1 vccd1 vccd1 y_i_1[3] sky130_fd_sc_hd__buf_2
Xoutput298 _10948_/X vssd1 vssd1 vccd1 vccd1 y_i_2[13] sky130_fd_sc_hd__buf_2
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07966_ _07966_/A vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__buf_6
XFILLER_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _15058_/Q _15091_/Q vssd1 vssd1 vccd1 vccd1 _09706_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07897_ _07897_/A vssd1 vssd1 vccd1 vccd1 _15319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_94_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15110_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _15303_/D sky130_fd_sc_hd__xor2_1
XFILLER_28_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _09786_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _15174_/D sky130_fd_sc_hd__xor2_1
XANTENNA__14187__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08518_ _08689_/A _08689_/B vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__xor2_1
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _15253_/D sky130_fd_sc_hd__xnor2_1
XFILLER_180_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08449_ _08600_/A _08599_/A vssd1 vssd1 vccd1 vccd1 _08458_/B sky130_fd_sc_hd__or2_1
XFILLER_211_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _11509_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__and3_1
XFILLER_23_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_952 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07416__A1 _07416_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ _15110_/Q _15209_/Q vssd1 vssd1 vccd1 vccd1 _10412_/C sky130_fd_sc_hd__and2b_1
XFILLER_136_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11391_ _11391_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11391_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_99_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input187_A x_r_3[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ _13712_/A _13712_/B _13713_/B vssd1 vssd1 vccd1 vccd1 _13131_/B sky130_fd_sc_hd__a21oi_2
X_10342_ _10469_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _15785_/D sky130_fd_sc_hd__xnor2_1
XFILLER_87_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _13061_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__and2_1
XFILLER_155_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10273_ _10273_/A _10279_/A vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_903 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14650__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _12148_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__nand2_1
XFILLER_2_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input48_A x_i_2[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13963_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13963_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15352_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15702_ _15761_/CLK _15702_/D _14777_/Y vssd1 vssd1 vccd1 vccd1 _15702_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12914_ _13677_/A _12986_/B vssd1 vssd1 vccd1 vccd1 _12914_/Y sky130_fd_sc_hd__nand2_1
X_13894_ _08793_/Y _13893_/B _08795_/B vssd1 vssd1 vccd1 vccd1 _13896_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13713__B _13713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15633_ _15773_/CLK _15633_/D _14705_/Y vssd1 vssd1 vccd1 vccd1 _15633_/Q sky130_fd_sc_hd__dfrtp_1
X_12845_ _12845_/A _12845_/B vssd1 vssd1 vccd1 vccd1 _12846_/B sky130_fd_sc_hd__nand2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14097__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15631__D _15631_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15564_ _15576_/CLK _15564_/D _14631_/Y vssd1 vssd1 vccd1 vccd1 _15564_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12777_/A _12777_/B _12777_/C vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__a21o_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07655__A1 input258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ _11727_/A vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__inv_2
X_14515_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14515_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _15511_/CLK _15495_/D _14558_/Y vssd1 vssd1 vccd1 vccd1 _15495_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_202_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11658_ _11658_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__nand2_1
X_14446_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _10609_/A _10609_/B _10609_/C vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__and3_1
XFILLER_174_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08604__B1 _08530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14377_/Y sky130_fd_sc_hd__inv_2
X_11589_ _11515_/Y _11587_/Y _11517_/B _11588_/Y vssd1 vssd1 vccd1 vccd1 _11607_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater619_A repeater620/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13328_ _13380_/A _13374_/C vssd1 vssd1 vccd1 vccd1 _13329_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08080__A1 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _13259_/A _13297_/A _13259_/C vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__or3_1
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14560__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12999__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater890_A input234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15806__D _15806_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _15357_/Q _07820_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__mux2_1
Xrepeater702 _07695_/S vssd1 vssd1 vccd1 vccd1 _07687_/S sky130_fd_sc_hd__buf_4
Xrepeater713 _15707_/Q vssd1 vssd1 vccd1 vccd1 output385/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater724 repeater725/X vssd1 vssd1 vccd1 vccd1 output351/A sky130_fd_sc_hd__buf_4
XFILLER_85_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater735 _15671_/Q vssd1 vssd1 vccd1 vccd1 output313/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater746 _15655_/Q vssd1 vssd1 vccd1 vccd1 repeater746/X sky130_fd_sc_hd__buf_2
X_07751_ _07751_/A vssd1 vssd1 vccd1 vccd1 _15391_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_92_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater757 _15644_/Q vssd1 vssd1 vccd1 vccd1 output285/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater768 _15630_/Q vssd1 vssd1 vccd1 vccd1 output526/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_76_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater779 _15618_/Q vssd1 vssd1 vccd1 vccd1 repeater779/X sky130_fd_sc_hd__buf_4
X_07682_ _07682_/A vssd1 vssd1 vccd1 vccd1 _15425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09421_ _15529_/Q _15513_/Q vssd1 vssd1 vccd1 vccd1 _09421_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07902__A _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07894__A1 _07894_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09352_ _09354_/C _09352_/B vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__and2_1
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08303_ _08283_/Y _08285_/Y _08287_/X _08289_/X _08302_/X vssd1 vssd1 vccd1 vccd1
+ _08303_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ _09283_/A _09283_/B vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__nor2_1
XFILLER_166_705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14735__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_30_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _15018_/Q vssd1 vssd1 vccd1 vccd1 _12312_/S sky130_fd_sc_hd__buf_4
XFILLER_147_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__B _15416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08452__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08096_ _08120_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__xnor2_2
XFILLER_161_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_45_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14470__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08374__A2 _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08998_ _13600_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _15106_/D sky130_fd_sc_hd__xor2_1
XFILLER_134_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07949_ _07949_/A vssd1 vssd1 vccd1 vccd1 _14987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_103_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10958_/A _11140_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09619_ _15444_/Q _15428_/Q vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__or2_1
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _14960_/Q _14894_/Q vssd1 vssd1 vccd1 vccd1 _10891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_203_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12630_ _12630_/A _12810_/A _12654_/A vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__and3_1
XFILLER_70_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input102_A x_i_6[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13252__C _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12561_ _15737_/Q _12219_/B _12560_/B vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14645__A _14661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ _11447_/X _11449_/A _11511_/Y vssd1 vssd1 vccd1 vccd1 _11530_/A sky130_fd_sc_hd__o21ai_1
XFILLER_8_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14300_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__buf_8
X_15280_ _15400_/CLK _15280_/D _14331_/Y vssd1 vssd1 vccd1 vccd1 _15280_/Q sky130_fd_sc_hd__dfrtp_1
X_12492_ _12262_/A _12491_/Y _12485_/A vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08643__A _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14231_/Y sky130_fd_sc_hd__inv_2
X_11443_ _12231_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__xnor2_1
XFILLER_137_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12165__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11374_ _15752_/Q _15030_/Q vssd1 vssd1 vccd1 vccd1 _11375_/C sky130_fd_sc_hd__and2_1
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _13113_/A _13113_/B vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__xnor2_1
X_10325_ _10317_/Y _10321_/B _10319_/B vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__o21ai_4
X_14093_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14093_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14380__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07693__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13101_/A _13044_/B vssd1 vssd1 vccd1 vccd1 _13046_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10256_ _10256_/A vssd1 vssd1 vccd1 vccd1 _15768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10187_ _10187_/A _10856_/A vssd1 vssd1 vccd1 vccd1 _15808_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__07573__A0 _15478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output321_A output321/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15133_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14995_ _15498_/CLK _14995_/D _14029_/Y vssd1 vssd1 vccd1 vccd1 _14995_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output419_A output419/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13946_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07876__A1 _07876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _13877_/A _13877_/B vssd1 vssd1 vccd1 vccd1 _15055_/D sky130_fd_sc_hd__xnor2_1
XFILLER_46_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater569_A repeater570/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _15732_/CLK _15616_/D _14687_/Y vssd1 vssd1 vccd1 vccd1 _15616_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _12717_/A _12717_/B _12827_/Y vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07628__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15547_ _15569_/CLK _15547_/D _14613_/Y vssd1 vssd1 vccd1 vccd1 _15547_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater736_A _15667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ _12759_/A _12687_/A vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__or2b_1
XANTENNA__14555__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15478_ _15761_/CLK _15478_/D _14540_/Y vssd1 vssd1 vccd1 vccd1 _15478_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14429_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09970_ _09970_/A _10009_/A vssd1 vssd1 vccd1 vccd1 _14970_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__14290__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ _08921_/A _08921_/B _08970_/A vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__and3_1
XFILLER_130_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08852_ _15461_/Q _08852_/B _08936_/B vssd1 vssd1 vccd1 vccd1 _08853_/B sky130_fd_sc_hd__and3_1
XANTENNA__10323__A _15126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07803_ _15365_/Q input227/X _07803_/S vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater532 _12221_/Y vssd1 vssd1 vccd1 vccd1 _15588_/D sky130_fd_sc_hd__clkbuf_2
X_08783_ _15339_/Q _15323_/Q vssd1 vssd1 vccd1 vccd1 _08783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater543 _11391_/Y vssd1 vssd1 vccd1 vccd1 output437/A sky130_fd_sc_hd__clkbuf_2
XFILLER_211_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15175_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater554 _11341_/Y vssd1 vssd1 vccd1 vccd1 output330/A sky130_fd_sc_hd__buf_4
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater565 _11087_/X vssd1 vssd1 vccd1 vccd1 repeater565/X sky130_fd_sc_hd__buf_2
X_07734_ _15399_/Q _07734_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater576 repeater577/X vssd1 vssd1 vccd1 vccd1 output364/A sky130_fd_sc_hd__buf_4
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater587 _11067_/Y vssd1 vssd1 vccd1 vccd1 repeater587/X sky130_fd_sc_hd__buf_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater598 _11056_/Y vssd1 vssd1 vccd1 vccd1 output275/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08728__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_836 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07665_ _15433_/Q _07665_/A1 _07697_/S vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _15412_/Q _15396_/Q vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07596_ _15467_/Q input79/X _07632_/S vssd1 vssd1 vccd1 vccd1 _07597_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _15410_/Q _15394_/Q vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__xnor2_4
XFILLER_34_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14465__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _09266_/A _09266_/B _09266_/C vssd1 vssd1 vccd1 vccd1 _09268_/A sky130_fd_sc_hd__and3_1
XFILLER_194_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_08217_ _11464_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__xor2_4
XFILLER_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09278__B _15381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _15572_/Q _15552_/Q vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__and2_1
XFILLER_14_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08148_ _15011_/Q vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__buf_6
XFILLER_162_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _08090_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08079_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12713__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _15138_/Q _15303_/Q vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__or2_1
XFILLER_106_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _14935_/Q _15001_/Q vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10041_ _15208_/Q _15109_/Q vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__or2_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _13798_/Y _13797_/B _13799_/X vssd1 vssd1 vccd1 vccd1 _13807_/A sky130_fd_sc_hd__a21o_1
XFILLER_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _12204_/A _12144_/A vssd1 vssd1 vccd1 vccd1 _11992_/Y sky130_fd_sc_hd__nor2_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14780_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _14901_/Q _14967_/Q vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__or2b_1
XANTENNA__07858__A1 input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13731_ _13838_/B _13731_/B vssd1 vssd1 vccd1 vccd1 _15701_/D sky130_fd_sc_hd__xor2_1
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08357__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10874_ _14956_/Q _10873_/Y _10869_/B vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13662_ _08757_/A _13809_/B _13813_/B _14972_/Q _13642_/X vssd1 vssd1 vccd1 vccd1
+ _13663_/B sky130_fd_sc_hd__a221o_1
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15588_/CLK _15401_/D _14459_/Y vssd1 vssd1 vccd1 vccd1 _15401_/Q sky130_fd_sc_hd__dfrtp_2
X_12613_ _12613_/A _12613_/B vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__nor2_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13593_ _15365_/Q _15349_/Q _13591_/B _13592_/X vssd1 vssd1 vccd1 vccd1 _13594_/B
+ sky130_fd_sc_hd__a31o_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14375__A _14379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ _12544_/A _12544_/B vssd1 vssd1 vccd1 vccd1 _15616_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__09469__A _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ _15782_/CLK _15332_/D _14386_/Y vssd1 vssd1 vccd1 vccd1 _15332_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12475_ _14949_/Q _12484_/B _12475_/C vssd1 vssd1 vccd1 vccd1 _12475_/Y sky130_fd_sc_hd__nand3_1
X_15263_ _15268_/CLK _15263_/D _14313_/Y vssd1 vssd1 vccd1 vccd1 _15263_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14214_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14214_/Y sky130_fd_sc_hd__inv_2
X_11426_ _11424_/A _11424_/B _11425_/X vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__a21oi_2
X_15194_ _15460_/CLK _15194_/D _14241_/Y vssd1 vssd1 vccd1 vccd1 _15194_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output271_A output271/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output369_A _11143_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14145_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14145_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11357_ _11357_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11357_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_4_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12623__A _15726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ _15123_/Q _15156_/Q vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14076_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14076_/Y sky130_fd_sc_hd__inv_2
X_11288_ _11287_/A _11287_/C _11287_/B vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__a21oi_1
XFILLER_141_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13027_ _13438_/A _13381_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__and3_1
X_10239_ _10239_/A _11406_/A _10239_/C vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__and3_1
XFILLER_117_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater686_A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_983 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14978_ _15774_/CLK _14978_/D _14011_/Y vssd1 vssd1 vccd1 vccd1 _14978_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13929_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07450_ _07450_/A vssd1 vssd1 vccd1 vccd1 _15539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07381_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07432_/S sky130_fd_sc_hd__buf_12
XFILLER_210_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14285__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _09120_/A _09258_/A vssd1 vssd1 vccd1 vccd1 _09254_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07598__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_360 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _09051_/A _09056_/A vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__or2_1
XFILLER_175_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10318__A _15125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08002_ _12238_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__xnor2_1
XFILLER_198_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13348__B _13746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _09953_/A _09953_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _09953_/X sky130_fd_sc_hd__and3_1
XFILLER_83_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08904_ _15456_/Q _15472_/Q vssd1 vssd1 vccd1 vccd1 _08906_/A sky130_fd_sc_hd__or2b_1
XFILLER_100_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09884_ _09975_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _15347_/Q _15331_/Q vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08766_/A _08766_/B _13877_/A vssd1 vssd1 vccd1 vccd1 _08768_/A sky130_fd_sc_hd__nor3_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07717_/A vssd1 vssd1 vccd1 vccd1 _15408_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _08529_/B _08697_/B vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__and2b_1
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07648_ _07648_/A vssd1 vssd1 vccd1 vccd1 _15442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07579_ _15475_/Q input72/X _07579_/S vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14195__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ _15407_/Q _15391_/Q vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__or2b_1
XFILLER_185_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10590_ _10590_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _14988_/D sky130_fd_sc_hd__xnor2_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09249_ _15502_/Q _15486_/Q vssd1 vssd1 vccd1 vccd1 _09250_/C sky130_fd_sc_hd__or2b_1
XFILLER_103_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ _12260_/A _12260_/B vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _11209_/X _11216_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__and2b_1
X_12191_ _12247_/A _12191_/B vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__xor2_1
XFILLER_108_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11142_ _10958_/B _11140_/B _11141_/Y vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12162__B _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11073_ _14932_/Q _14998_/Q vssd1 vssd1 vccd1 vccd1 _11077_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput110 x_i_6[5] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput121 x_i_7[15] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14901_ _15732_/CLK _14901_/D _13930_/Y vssd1 vssd1 vccd1 vccd1 _14901_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input30_A x_i_1[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput132 x_r_0[10] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10024_ _10020_/A _10017_/Y _10019_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__o21ai_2
Xinput143 x_r_0[6] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__clkbuf_2
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput154 x_r_1[1] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput165 x_r_2[11] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__clkbuf_1
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 x_r_2[7] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_hd__clkbuf_2
Xinput187 x_r_3[2] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14832_/Y sky130_fd_sc_hd__inv_2
Xinput198 x_r_4[12] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13077__A1 _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14763_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14763_/Y sky130_fd_sc_hd__inv_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _12029_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11977_/B sky130_fd_sc_hd__xnor2_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13714_ _13715_/A _13715_/B vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__or2_1
XFILLER_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10926_ _10924_/X _10931_/B vssd1 vssd1 vccd1 vccd1 _10927_/A sky130_fd_sc_hd__and2b_2
XANTENNA__07700__A0 _15416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14694_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14694_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10857_ _15809_/Q _14955_/Q vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__or2b_1
XFILLER_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13645_ _13645_/A _13645_/B vssd1 vssd1 vccd1 vccd1 _13646_/C sky130_fd_sc_hd__and2_1
XFILLER_204_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11522__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10788_ _10787_/A _10787_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _10795_/A sky130_fd_sc_hd__a21o_1
X_13576_ _15769_/Q _13576_/B vssd1 vssd1 vccd1 vccd1 _13576_/X sky130_fd_sc_hd__and2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_680 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output486_A output486/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _15575_/CLK _15315_/D _14368_/Y vssd1 vssd1 vccd1 vccd1 _15315_/Q sky130_fd_sc_hd__dfrtp_1
X_12527_ _12527_/A _12527_/B vssd1 vssd1 vccd1 vccd1 _12527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14833__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13001__A1 _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15246_ _15249_/CLK _15246_/D _14295_/Y vssd1 vssd1 vccd1 vccd1 _15246_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12458_ _12458_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11409_ _15078_/Q _15243_/Q _11408_/B vssd1 vssd1 vccd1 vccd1 _11411_/C sky130_fd_sc_hd__a21o_1
XFILLER_99_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12389_ _14942_/Q _12391_/C _12389_/C vssd1 vssd1 vccd1 vccd1 _12398_/A sky130_fd_sc_hd__and3_1
XFILLER_172_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ _15663_/CLK _15177_/D _14222_/Y vssd1 vssd1 vccd1 vccd1 _15177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14128_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14059_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_80_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater970_A repeater971/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13184__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08620_ _08573_/A _08573_/B _08615_/A vssd1 vssd1 vccd1 vccd1 _08621_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _08551_/A _08577_/A vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__or2_1
X_07502_ _15513_/Q input29/X _07536_/S vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08482_ _14909_/Q vssd1 vssd1 vccd1 vccd1 _12871_/A sky130_fd_sc_hd__buf_6
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07433_ _07433_/A vssd1 vssd1 vccd1 vccd1 _15547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07910__A _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _09243_/A _09103_/B vssd1 vssd1 vccd1 vccd1 _15226_/D sky130_fd_sc_hd__xnor2_1
XFILLER_202_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14743__A _14751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09034_/A vssd1 vssd1 vccd1 vccd1 _15112_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13679__B1_N _12910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _15196_/Q _15229_/Q vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__or2b_1
XANTENNA__07791__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09572__A _15437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09867_ _15186_/Q _15219_/Q vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__or2b_1
XFILLER_112_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15724__D _15724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13094__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08818_/A _08818_/B _13901_/A vssd1 vssd1 vccd1 vccd1 _08818_/X sky130_fd_sc_hd__and3_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09798_ _15439_/Q _15423_/Q vssd1 vssd1 vccd1 vccd1 _09799_/C sky130_fd_sc_hd__and2_1
XFILLER_133_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _08707_/Y _08748_/Y _08710_/X _08748_/B vssd1 vssd1 vccd1 vccd1 _08750_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _12178_/A _12055_/A _12038_/B vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__and3_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _15183_/Q _15282_/Q vssd1 vssd1 vccd1 vccd1 _10712_/B sky130_fd_sc_hd__and2b_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11691_ _12204_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _11692_/C sky130_fd_sc_hd__xor2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10642_ _10642_/A _10642_/B vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__nand2_2
X_13430_ _13431_/B _14920_/Q vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__nor2b_1
XFILLER_9_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13361_ _13361_/A _13361_/B vssd1 vssd1 vccd1 vccd1 _13362_/C sky130_fd_sc_hd__or2_1
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10573_ _10572_/A _10572_/B _10619_/A vssd1 vssd1 vccd1 vccd1 _10577_/B sky130_fd_sc_hd__a21o_1
XFILLER_194_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14653__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15100_ _15375_/CLK _15100_/D _14141_/Y vssd1 vssd1 vccd1 vccd1 _15100_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_194_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ _12246_/X _12245_/Y _12312_/S vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__mux2_2
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13292_ _13712_/A _13712_/B _13713_/B _13063_/A vssd1 vssd1 vccd1 vccd1 _13292_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_166_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input78_A x_i_4[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12243_ _12243_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12262_/A sky130_fd_sc_hd__xnor2_2
X_15031_ _15483_/CLK _15031_/D _14068_/Y vssd1 vssd1 vccd1 vccd1 _15031_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_839 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12174_ _12175_/A _12175_/B _12175_/C vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__a21o_1
XFILLER_174_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11125_ _11125_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _11125_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11056_ _11327_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11056_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_7_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15634__D _15634_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _15200_/Q _15233_/Q vssd1 vssd1 vccd1 vccd1 _10007_/Y sky130_fd_sc_hd__nand2_1
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1016 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14815_/Y sky130_fd_sc_hd__inv_2
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15795_/CLK _15795_/D _14875_/Y vssd1 vssd1 vccd1 vccd1 _15795_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14828__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14750_/A vssd1 vssd1 vccd1 vccd1 _14746_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ _12238_/A _12231_/A _11956_/X vssd1 vssd1 vccd1 vccd1 _11959_/B sky130_fd_sc_hd__a21o_1
XFILLER_205_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10909_ _14895_/Q _14961_/Q vssd1 vssd1 vccd1 vccd1 _10910_/C sky130_fd_sc_hd__or2b_1
XANTENNA_repeater551_A _11140_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14677_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14677_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11889_ _11890_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__or2_1
XANTENNA_repeater649_A _07971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1000 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08229__A1 _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13628_ _13628_/A _13628_/B vssd1 vssd1 vccd1 vccd1 _15100_/D sky130_fd_sc_hd__xnor2_1
XFILLER_193_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater816_A _14862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ _13561_/A _13560_/B _13561_/B _13560_/A vssd1 vssd1 vccd1 vccd1 _13564_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_173_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14563__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07876__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13179__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput403 output403/A vssd1 vssd1 vccd1 vccd1 y_r_0[16] sky130_fd_sc_hd__buf_2
X_15229_ _15501_/CLK _15229_/D _14277_/Y vssd1 vssd1 vccd1 vccd1 _15229_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput414 output414/A vssd1 vssd1 vccd1 vccd1 y_r_1[10] sky130_fd_sc_hd__buf_2
XFILLER_201_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput425 output425/A vssd1 vssd1 vccd1 vccd1 y_r_1[5] sky130_fd_sc_hd__buf_2
Xoutput436 _11388_/Y vssd1 vssd1 vccd1 vccd1 y_r_2[15] sky130_fd_sc_hd__buf_2
Xoutput447 output447/A vssd1 vssd1 vccd1 vccd1 y_r_3[0] sky130_fd_sc_hd__buf_2
XFILLER_114_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput458 output458/A vssd1 vssd1 vccd1 vccd1 y_r_3[4] sky130_fd_sc_hd__buf_2
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput469 output469/A vssd1 vssd1 vccd1 vccd1 y_r_4[14] sky130_fd_sc_hd__buf_2
XFILLER_99_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07982_ _11678_/A _11584_/A _07995_/A vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__and3_1
XFILLER_99_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09721_ _09719_/Y _09721_/B vssd1 vssd1 vccd1 vccd1 _09840_/A sky130_fd_sc_hd__and2b_1
XFILLER_171_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09652_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09654_/B sky130_fd_sc_hd__and2_1
XFILLER_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08603_ _12810_/A _08603_/B vssd1 vssd1 vccd1 vccd1 _08603_/X sky130_fd_sc_hd__or2_1
X_09583_ _09791_/A _09577_/B _09582_/X vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14738__A _14741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _08728_/A _12688_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08550_/A sky130_fd_sc_hd__and3_2
XFILLER_42_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08465_ _08466_/B _08451_/A _08451_/B _08589_/A _08589_/B vssd1 vssd1 vccd1 vccd1
+ _08587_/B sky130_fd_sc_hd__a32o_1
XFILLER_208_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07416_ _15555_/Q _07416_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ _08396_/A _12654_/A _08396_/C vssd1 vssd1 vccd1 vccd1 _08441_/A sky130_fd_sc_hd__and3_1
XFILLER_195_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14473__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08471__A _14905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15719__D _15719_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _13607_/A _09012_/B _09016_/X vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08943__A2 _15448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09919_ _09918_/A _09918_/C _09985_/A vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12930_ _12930_/A _12930_/B vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input132_A x_r_0[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12957_/A _12667_/C _13046_/A vssd1 vssd1 vccd1 vccd1 _12862_/B sky130_fd_sc_hd__mux2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14648__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_901 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14600_/Y sky130_fd_sc_hd__inv_2
X_11812_ _11587_/Y _11766_/A _11767_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11814_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15648_/CLK _15580_/D _14649_/Y vssd1 vssd1 vccd1 vccd1 _15580_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08646__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ _14920_/Q _12791_/B _12791_/C vssd1 vssd1 vccd1 vccd1 _12793_/B sky130_fd_sc_hd__a21oi_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14531_/Y sky130_fd_sc_hd__inv_2
X_11743_ _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08365__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14462_/Y sky130_fd_sc_hd__inv_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11603_/A _11602_/B _11602_/A vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__o21bai_1
XFILLER_202_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13413_ _13356_/A _13356_/B _13361_/A vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__a21o_1
X_10625_ _10625_/A _10625_/B vssd1 vssd1 vccd1 vccd1 _15002_/D sky130_fd_sc_hd__xnor2_1
XFILLER_168_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14393_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14383__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11800__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13345_/B sky130_fd_sc_hd__xnor2_2
X_10556_ _15295_/Q _15262_/Q vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__or2b_1
XFILLER_154_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _15285_/Q _15252_/Q vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__or2b_1
X_13275_ _13274_/A _13274_/B _13274_/C vssd1 vssd1 vccd1 vccd1 _13316_/C sky130_fd_sc_hd__a21o_1
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15014_ _15435_/CLK _15014_/D _14050_/Y vssd1 vssd1 vccd1 vccd1 _15014_/Q sky130_fd_sc_hd__dfrtp_1
X_12226_ _12556_/B _12560_/A vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__or2_1
XFILLER_170_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output351_A output351/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output449_A _15605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ _12156_/A _12156_/B _12556_/B vssd1 vssd1 vccd1 vccd1 _12220_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ _10864_/Y _11107_/B _10866_/B vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__o21ai_2
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12089_/C sky130_fd_sc_hd__xnor2_1
XFILLER_110_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater906 input213/X vssd1 vssd1 vccd1 vccd1 _07716_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater917 input193/X vssd1 vssd1 vccd1 vccd1 _07689_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater928 input177/X vssd1 vssd1 vccd1 vccd1 _07820_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater939 input161/X vssd1 vssd1 vccd1 vccd1 _07755_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11039_ _11039_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08698__A1 _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater766_A _15633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14558__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15778_ _15791_/CLK _15778_/D _14857_/Y vssd1 vssd1 vccd1 vccd1 _15778_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14729_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14729_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater933_A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08250_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08257_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08181_ _11687_/A _11491_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08189_/A sky130_fd_sc_hd__and3_1
XFILLER_158_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14293__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A1 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput266 _11100_/X vssd1 vssd1 vccd1 vccd1 y_i_0[15] sky130_fd_sc_hd__buf_2
XFILLER_102_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput277 output277/A vssd1 vssd1 vccd1 vccd1 y_i_1[0] sky130_fd_sc_hd__buf_2
XFILLER_160_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput288 output288/A vssd1 vssd1 vccd1 vccd1 y_i_1[4] sky130_fd_sc_hd__buf_2
XFILLER_59_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput299 _10952_/Y vssd1 vssd1 vccd1 vccd1 y_i_2[14] sky130_fd_sc_hd__buf_2
XFILLER_173_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07965_ _11353_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__and2_1
XANTENNA__15274__D _15274_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ _15058_/Q _15091_/Q vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__or2_1
X_07896_ _15319_/Q _07896_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09635_ _09634_/Y _15543_/Q _09633_/B vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14468__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09566_ _09783_/A _09561_/B _09565_/X vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13434__A1 _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08517_ _13438_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08689_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09497_ _15525_/Q _15509_/Q _09495_/B _09496_/X vssd1 vssd1 vccd1 vccd1 _09498_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09231__A_N _15497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08448_ _13012_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08599_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ _15042_/Q vssd1 vssd1 vccd1 vccd1 _12945_/A sky130_fd_sc_hd__buf_6
XFILLER_196_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10410_ _10410_/A _10412_/B vssd1 vssd1 vccd1 vccd1 _14946_/D sky130_fd_sc_hd__nor2_1
XFILLER_139_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11390_ _11243_/B _11388_/B _11389_/Y vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__o21ai_1
XFILLER_165_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _13061_/A _13100_/B _13062_/B vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__and3_1
X_10272_ _15247_/Q _15082_/Q vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__or2b_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _12011_/A _12011_/B _12009_/Y vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__or3b_1
XFILLER_155_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13962_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15701_ _15706_/CLK _15701_/D _14776_/Y vssd1 vssd1 vccd1 vccd1 _15701_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12913_ _13021_/B _12913_/B vssd1 vssd1 vccd1 vccd1 _12986_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14378__A _14379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ _13893_/A _13893_/B vssd1 vssd1 vccd1 vccd1 _15061_/D sky130_fd_sc_hd__xor2_1
XFILLER_73_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15632_ _15708_/CLK _15632_/D _14704_/Y vssd1 vssd1 vccd1 vccd1 _15632_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12844_ _12699_/Y _13528_/B _13535_/B _12843_/A _12700_/X vssd1 vssd1 vccd1 vccd1
+ _12845_/B sky130_fd_sc_hd__o221ai_2
XFILLER_64_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08376__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__B _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15563_/CLK _15563_/D _14630_/Y vssd1 vssd1 vccd1 vccd1 _15563_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12775_/A vssd1 vssd1 vccd1 vccd1 _12777_/C sky130_fd_sc_hd__inv_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14514_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11723_/A _11724_/Y _11725_/X vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__a21o_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15664_/CLK _15494_/D _14557_/Y vssd1 vssd1 vccd1 vccd1 _15494_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output399_A _10782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14445_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14445_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11680_/A sky130_fd_sc_hd__or2_1
XANTENNA__08604__A1 _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ _10609_/A _10609_/C _10609_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__a21oi_1
XFILLER_155_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14376_ _14376_/A vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__inv_2
X_11588_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11588_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13327_ _14920_/Q _13327_/B vssd1 vssd1 vccd1 vccd1 _13374_/C sky130_fd_sc_hd__nor2_1
XFILLER_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10146__A _15310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ _15260_/Q _15293_/Q vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__or2_1
XFILLER_182_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14841__A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09935__A _09935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ _13258_/A _13258_/B vssd1 vssd1 vccd1 vccd1 _13259_/C sky130_fd_sc_hd__or2_1
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _12209_/A _12209_/B vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__or2_1
XFILLER_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _13189_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13190_/B sky130_fd_sc_hd__and2_1
XFILLER_9_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater883_A input242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater703 _07644_/S vssd1 vssd1 vccd1 vccd1 _07640_/S sky130_fd_sc_hd__buf_6
Xrepeater714 _15705_/Q vssd1 vssd1 vccd1 vccd1 output383/A sky130_fd_sc_hd__buf_4
XANTENNA__07591__A1 _07591_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater725 _15691_/Q vssd1 vssd1 vccd1 vccd1 repeater725/X sky130_fd_sc_hd__buf_2
XFILLER_78_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater736 _15667_/Q vssd1 vssd1 vccd1 vccd1 output325/A sky130_fd_sc_hd__clkbuf_2
X_07750_ _15391_/Q _07750_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07751_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater747 repeater748/X vssd1 vssd1 vccd1 vccd1 output279/A sky130_fd_sc_hd__buf_4
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater758 _15643_/Q vssd1 vssd1 vccd1 vccd1 output277/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater769 _15629_/Q vssd1 vssd1 vccd1 vccd1 output525/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07681_ _15425_/Q input182/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14288__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _09501_/A _09420_/B vssd1 vssd1 vccd1 vccd1 _15270_/D sky130_fd_sc_hd__xor2_1
XANTENNA__07902__B _15317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _15397_/Q _09351_/B _09351_/C vssd1 vssd1 vccd1 vccd1 _09352_/B sky130_fd_sc_hd__nand3_1
XFILLER_178_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08302_ _08291_/Y _08292_/Y _08283_/Y _08285_/Y _08301_/X vssd1 vssd1 vccd1 vccd1
+ _08302_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13920__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _15399_/Q _15383_/Q vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08233_ _08220_/Y _08232_/A _08230_/X _08243_/B _08243_/A vssd1 vssd1 vccd1 vccd1
+ _08235_/B sky130_fd_sc_hd__a32o_1
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11440__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _12254_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _08120_/B _08120_/C vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14751__A _14751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_1_0_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08997_ _13597_/A _08992_/B _08996_/X vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07948_ _10590_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__and2_1
XFILLER_69_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14198__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07879_ _07879_/A vssd1 vssd1 vccd1 vccd1 _15328_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15732__D _15732_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_826 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _15444_/Q _15428_/Q vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ _11113_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ _15431_/Q vssd1 vssd1 vccd1 vccd1 _09549_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__C1 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _12560_/A _12560_/B vssd1 vssd1 vccd1 vccd1 _15621_/D sky130_fd_sc_hd__xor2_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08924__A _15475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11511_ _08010_/Y _11584_/A _11445_/B _11678_/A _11876_/A vssd1 vssd1 vccd1 vccd1
+ _11511_/Y sky130_fd_sc_hd__o2111ai_1
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _12491_/A vssd1 vssd1 vccd1 vccd1 _12491_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08643__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14230_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14230_/Y sky130_fd_sc_hd__inv_2
X_11442_ _11442_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11519_/B sky130_fd_sc_hd__xnor2_1
XFILLER_165_761 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14161_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14161_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ _11373_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11373_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14661__A _14661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ _10324_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__nand2_2
XANTENNA_input60_A x_i_3[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13162_/B _13112_/B vssd1 vssd1 vccd1 vccd1 _13113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_153_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09755__A _09755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14092_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14092_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12146__A1 _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13043_ _12965_/A _12965_/B _13042_/X vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__o21ai_1
X_10255_ _10253_/X _10260_/B vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10186_ _15151_/Q _15316_/Q vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__xnor2_2
XFILLER_67_918 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07573__A1 _07573_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14994_ _15027_/CLK _14994_/D _14028_/Y vssd1 vssd1 vccd1 vccd1 _14994_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13945_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13945_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output314_A output314/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13876_ _15333_/Q _15317_/Q _13874_/B _13875_/X vssd1 vssd1 vccd1 vccd1 _13877_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15615_ _15689_/CLK _15615_/D _14686_/Y vssd1 vssd1 vccd1 vccd1 _15615_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_201_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12827_ _12827_/A _12827_/B vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14836__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ _15553_/CLK _15546_/D _14612_/Y vssd1 vssd1 vccd1 vccd1 _15546_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__xnor2_2
XFILLER_163_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _11709_/A _11709_/B _11709_/C vssd1 vssd1 vccd1 vccd1 _11710_/B sky130_fd_sc_hd__and3_1
XFILLER_202_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater631_A _10733_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15477_ _15477_/CLK _15477_/D _14539_/Y vssd1 vssd1 vccd1 vccd1 _15477_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12689_ _12690_/A _12690_/B _12690_/C vssd1 vssd1 vccd1 vccd1 _12691_/A sky130_fd_sc_hd__a21oi_1
XFILLER_175_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14428_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14428_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14359_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14359_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14571__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07884__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08920_ _08920_/A _08925_/A vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__or2_1
XFILLER_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08851_ _15461_/Q _08852_/B _08936_/B vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07802_ _07802_/A vssd1 vssd1 vccd1 vccd1 _15366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater533 _13450_/X vssd1 vssd1 vccd1 vccd1 _15638_/D sky130_fd_sc_hd__clkbuf_2
X_08782_ _13885_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _15074_/D sky130_fd_sc_hd__xor2_1
XFILLER_85_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater544 _11232_/X vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__buf_2
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater555 repeater556/X vssd1 vssd1 vccd1 vccd1 output466/A sky130_fd_sc_hd__buf_6
X_07733_ _07733_/A vssd1 vssd1 vccd1 vccd1 _15400_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater566 _10933_/X vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__buf_4
Xrepeater577 _11129_/Y vssd1 vssd1 vccd1 vccd1 repeater577/X sky130_fd_sc_hd__buf_2
XFILLER_37_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater588 _10773_/X vssd1 vssd1 vccd1 vccd1 output398/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08728__B _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater599 _10897_/Y vssd1 vssd1 vccd1 vccd1 output307/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07664_ _07664_/A vssd1 vssd1 vccd1 vccd1 _15434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ _09403_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _15150_/D sky130_fd_sc_hd__xnor2_1
XFILLER_197_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _07595_/A vssd1 vssd1 vccd1 vccd1 _15468_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14746__A _14750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09334_ _09332_/A _09390_/B _09333_/X vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__a21oi_4
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10993__B _15275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09265_ _09265_/A _09265_/B vssd1 vssd1 vccd1 vccd1 _09266_/C sky130_fd_sc_hd__nand2_1
XFILLER_194_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _08292_/B _08263_/B _08215_/Y vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09196_ _09196_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _15295_/D sky130_fd_sc_hd__xor2_1
XFILLER_181_506 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ _11832_/A _11687_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_1083 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08078_ _08090_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__xor2_1
XFILLER_84_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_786 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12713__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13876__A1 _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _10400_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _14976_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07555__A1 _07555_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11991_ _11991_/A _12088_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__and3_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _13721_/A _13832_/B _13729_/Y vssd1 vssd1 vccd1 vccd1 _13731_/B sky130_fd_sc_hd__o21a_1
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input212_A x_r_5[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ _14967_/Q _14901_/Q vssd1 vssd1 vccd1 vccd1 _10944_/A sky130_fd_sc_hd__or2b_1
XFILLER_17_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _14972_/Q _13813_/B vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__or2_1
X_10873_ _14890_/Q vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14656__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ _15400_/CLK _15400_/D _14458_/Y vssd1 vssd1 vccd1 vccd1 _15400_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12504_/B _14951_/Q vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__and2b_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13592_ _15366_/Q _15350_/Q vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__and2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15782_/CLK _15331_/D _14385_/Y vssd1 vssd1 vccd1 vccd1 _15331_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12543_/A _12543_/B vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__nand2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11080__A _11080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15262_ _15268_/CLK _15262_/D _14312_/Y vssd1 vssd1 vccd1 vccd1 _15262_/Q sky130_fd_sc_hd__dfrtp_1
X_12474_ _12604_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _15654_/D sky130_fd_sc_hd__xnor2_1
XFILLER_138_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_91_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14213_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _15083_/Q _15248_/Q vssd1 vssd1 vccd1 vccd1 _11425_/X sky130_fd_sc_hd__and2_1
XANTENNA__14391__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15193_ _15202_/CLK _15193_/D _14238_/Y vssd1 vssd1 vccd1 vccd1 _15193_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12904__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10145__B_N _15310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14144_/Y sky130_fd_sc_hd__inv_2
X_11356_ _11150_/Y _11355_/B _11152_/B vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__o21ai_4
XFILLER_113_606 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15637__D _15637_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10307_ _15123_/Q _15156_/Q vssd1 vssd1 vccd1 vccd1 _10307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14075_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14075_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11287_ _11287_/A _11287_/B _11287_/C vssd1 vssd1 vccd1 vccd1 _11289_/A sky130_fd_sc_hd__and3_1
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13026_ _13491_/S _13390_/A vssd1 vssd1 vccd1 vccd1 _13027_/C sky130_fd_sc_hd__xor2_1
X_10238_ _15241_/Q _15076_/Q vssd1 vssd1 vccd1 vccd1 _10239_/C sky130_fd_sc_hd__or2b_1
XANTENNA_output431_A output431/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_704 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output529_A output529/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _10168_/A _10168_/B _10850_/A vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14977_ _15249_/CLK _14977_/D _14010_/Y vssd1 vssd1 vccd1 vccd1 _14977_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater679_A _14526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13928_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13928_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13859_ _13859_/A _13859_/B vssd1 vssd1 vccd1 vccd1 _13860_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12785__S _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater846_A repeater847/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14566__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07380_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__buf_6
XFILLER_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15529_ _15532_/CLK _15529_/D _14594_/Y vssd1 vssd1 vccd1 vccd1 _15529_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_203_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09050_ _15378_/Q _15362_/Q vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__and2b_1
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_59_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ _08001_/A _08009_/C vssd1 vssd1 vccd1 vccd1 _08015_/B sky130_fd_sc_hd__xnor2_1
XFILLER_175_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07785__A1 _07785_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ _09952_/A _09958_/A vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _08903_/A vssd1 vssd1 vccd1 vccd1 _15211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_117_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09883_ _09975_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _14957_/D sky130_fd_sc_hd__xor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _15082_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08765_ _15335_/Q _15319_/Q vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__15282__D _15282_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07716_ _15408_/Q _07716_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__mux2_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _12662_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__xnor2_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07647_ _15442_/Q _07647_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14476__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08474__A _14906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ _07578_/A vssd1 vssd1 vccd1 vccd1 _15476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12708__B _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09317_ _15391_/Q _15407_/Q vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__or2b_1
XFILLER_16_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09248_ _09248_/A vssd1 vssd1 vccd1 vccd1 _15243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12349__A1 _12332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_09179_ _15570_/Q _15550_/Q vssd1 vssd1 vccd1 vccd1 _09188_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11210_ _11209_/A _11209_/B _11372_/B vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__a21o_1
X_12190_ _12190_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12191_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11141_ _14969_/Q _14903_/Q vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input162_A x_r_1[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11072_ _11072_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__nand2_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 x_i_6[10] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07528__A1 _07528_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12521__A1 _12332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput111 x_i_6[6] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_2
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14900_ _15133_/CLK _14900_/D _13929_/Y vssd1 vssd1 vccd1 vccd1 _14900_/Q sky130_fd_sc_hd__dfrtp_1
Xinput122 x_i_7[1] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__nand2_2
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 x_r_0[11] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput144 x_r_0[7] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_2
Xinput155 x_r_1[2] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 x_r_2[12] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput177 x_r_2[8] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__clkbuf_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input23_A x_i_1[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14831_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13077__A2 _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput188 x_r_3[3] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__clkbuf_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput199 x_r_4[13] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_2
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14762_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11974_ _11894_/A _11894_/B _11891_/A vssd1 vssd1 vccd1 vccd1 _11975_/B sky130_fd_sc_hd__o21ai_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13713_/A _13713_/B vssd1 vssd1 vccd1 vccd1 _13715_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_976 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _10924_/A _10924_/B _11124_/B vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__a21o_1
X_14693_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14693_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A1 _07700_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14386__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11803__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ _14972_/Q vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__inv_2
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10856_ _10856_/A _10856_/B vssd1 vssd1 vccd1 vccd1 _14920_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__08384__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11522__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13575_ _15769_/Q _13576_/B vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__or2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10787_ _10787_/A _10787_/B _11294_/A vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__and3_1
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15576_/CLK _15314_/D _14367_/Y vssd1 vssd1 vccd1 vccd1 _15314_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12526_ _15727_/Q vssd1 vssd1 vccd1 vccd1 _12527_/A sky130_fd_sc_hd__inv_2
XFILLER_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output381_A output381/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output479_A output479/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15245_ _15764_/CLK _15245_/D _14294_/Y vssd1 vssd1 vccd1 vccd1 _15245_/Q sky130_fd_sc_hd__dfrtp_1
X_12457_ _12456_/B _12456_/C _12456_/D _12456_/A vssd1 vssd1 vccd1 vccd1 _12468_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11408_ _11408_/A _11408_/B vssd1 vssd1 vccd1 vccd1 _15735_/D sky130_fd_sc_hd__xnor2_2
X_15176_ _15663_/CLK _15176_/D _14221_/Y vssd1 vssd1 vccd1 vccd1 _15176_/Q sky130_fd_sc_hd__dfrtp_1
X_12388_ _12388_/A _12398_/B vssd1 vssd1 vccd1 vccd1 _15647_/D sky130_fd_sc_hd__nor2_1
XFILLER_126_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07767__A1 input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14127_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14127_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11339_ _11339_/A _11339_/B _11339_/C vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__and3_1
XFILLER_193_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09508__A2 _15514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14058_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14058_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater796_A repeater797/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13009_ _13008_/A _13008_/B _13008_/C vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__a21o_1
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08559__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _08550_/A _08550_/B vssd1 vssd1 vccd1 vccd1 _08577_/A sky130_fd_sc_hd__xnor2_4
XFILLER_78_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07501_ _07501_/A vssd1 vssd1 vccd1 vccd1 _15514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ _12803_/A _12688_/A vssd1 vssd1 vccd1 vccd1 _08484_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14296__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07432_ _15547_/Q _07432_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11098__A_N _15002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07910__B _15349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07402__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ _09095_/Y _09100_/B _09097_/B vssd1 vssd1 vccd1 vccd1 _09103_/B sky130_fd_sc_hd__o21ai_1
XFILLER_202_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ _09031_/X _09038_/B vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10460__B_N _15126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_580 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_274 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09935_ _09935_/A vssd1 vssd1 vccd1 vccd1 _14964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09866_ _15219_/Q _15186_/Q vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__or2b_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _08817_/A _08825_/A vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09797_ _09797_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _15162_/D sky130_fd_sc_hd__nor2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08748_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08748_/Y sky130_fd_sc_hd__nand2_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__B _13822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__xnor2_1
XFILLER_96_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15740__D _15740_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10710_ _15282_/Q _15183_/Q vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__and2b_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11468_/Y _11626_/A _11627_/B _11627_/A vssd1 vssd1 vccd1 vccd1 _11705_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ _15270_/Q _15171_/Q vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ _13360_/A _13360_/B vssd1 vssd1 vccd1 vccd1 _13361_/B sky130_fd_sc_hd__and2_1
XFILLER_10_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10572_ _10572_/A _10572_/B _10619_/A vssd1 vssd1 vccd1 vccd1 _10572_/X sky130_fd_sc_hd__and3_1
XFILLER_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ _12287_/B _12289_/B _12310_/Y vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__o21a_2
XFILLER_5_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13291_ _13703_/B _13715_/A vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__and2_1
XFILLER_177_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15030_ _15498_/CLK _15030_/D _14067_/Y vssd1 vssd1 vccd1 vccd1 _15030_/Q sky130_fd_sc_hd__dfrtp_1
X_12242_ _12182_/B _12185_/B _12180_/Y vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ _12236_/B _12173_/B vssd1 vssd1 vccd1 vccd1 _12175_/C sky130_fd_sc_hd__or2_1
XFILLER_64_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _11124_/A _11124_/B _11124_/C vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__and3_1
XFILLER_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11049_/A _11051_/B _11049_/B vssd1 vssd1 vccd1 vccd1 _11056_/B sky130_fd_sc_hd__a21boi_2
XFILLER_209_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10702__A _15280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _14936_/D sky130_fd_sc_hd__xnor2_1
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14814_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14814_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15794_ _15795_/CLK _15794_/D _14874_/Y vssd1 vssd1 vccd1 vccd1 _15794_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14745_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14745_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11957_ _11957_/A _11956_/X vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__or2b_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15650__D _15650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11481__A1 _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _10906_/Y _10908_/B vssd1 vssd1 vccd1 vccd1 _11119_/A sky130_fd_sc_hd__and2b_2
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14676_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14676_/Y sky130_fd_sc_hd__inv_2
X_11888_ _11955_/A _11954_/A vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__xor2_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09003__A _15371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13627_ _13625_/A _13625_/B _13626_/X vssd1 vssd1 vccd1 vccd1 _13628_/B sky130_fd_sc_hd__a21o_1
X_10839_ _10839_/A _10839_/B _10839_/C vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__and3_1
XFILLER_34_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14844__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13558_ _15765_/Q _13558_/B vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12509_ _12509_/A vssd1 vssd1 vccd1 vccd1 _15657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater711_A _07434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13489_ _13463_/A _13463_/B _13464_/A vssd1 vssd1 vccd1 vccd1 _13490_/B sky130_fd_sc_hd__o21a_1
XANTENNA_repeater809_A _15578_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08561__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15228_ _15501_/CLK _15228_/D _14276_/Y vssd1 vssd1 vccd1 vccd1 _15228_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13179__B _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput404 output404/A vssd1 vssd1 vccd1 vccd1 y_r_0[1] sky130_fd_sc_hd__buf_2
Xoutput415 output415/A vssd1 vssd1 vccd1 vccd1 y_r_1[11] sky130_fd_sc_hd__buf_2
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput426 output426/A vssd1 vssd1 vccd1 vccd1 y_r_1[6] sky130_fd_sc_hd__buf_2
Xoutput437 output437/A vssd1 vssd1 vccd1 vccd1 y_r_2[16] sky130_fd_sc_hd__buf_2
Xoutput448 output448/A vssd1 vssd1 vccd1 vccd1 y_r_3[10] sky130_fd_sc_hd__buf_2
X_15159_ _15434_/CLK _15159_/D _14203_/Y vssd1 vssd1 vccd1 vccd1 _15159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput459 _15599_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[5] sky130_fd_sc_hd__buf_2
XFILLER_141_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07892__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07981_ _11797_/A _11658_/A vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__xor2_1
XFILLER_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09720_ _15061_/Q _15094_/Q vssd1 vssd1 vccd1 vccd1 _09721_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09651_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _15308_/D sky130_fd_sc_hd__xor2_1
XFILLER_55_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08602_ _12921_/A vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__inv_2
XANTENNA__13923__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ _15437_/Q _15421_/Q vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__and2b_1
X_08533_ _13220_/A vssd1 vssd1 vccd1 vccd1 _13030_/C sky130_fd_sc_hd__inv_2
XFILLER_70_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11443__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08464_ _08464_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08589_/B sky130_fd_sc_hd__xnor2_1
XFILLER_196_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07415_ _07415_/A vssd1 vssd1 vccd1 vccd1 _15556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08395_ _13273_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__xnor2_1
XFILLER_177_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14754__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11883__A_N _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09010__A_N _15371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ _15372_/Q _15356_/Q vssd1 vssd1 vccd1 vccd1 _09016_/X sky130_fd_sc_hd__and2b_1
XFILLER_12_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15735__D _15735_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09918_ _09918_/A _09985_/A _09918_/C vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__and3_1
XFILLER_24_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09849_ _09848_/B _09848_/C _09848_/A vssd1 vssd1 vccd1 vccd1 _09852_/C sky130_fd_sc_hd__a21o_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12860_ _13145_/A vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__inv_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A x_i_7[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A _11811_/B vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__xnor2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _14920_/Q _12791_/B _12791_/C vssd1 vssd1 vccd1 vccd1 _12793_/A sky130_fd_sc_hd__and3_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08646__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14530_/Y sky130_fd_sc_hd__inv_2
X_11742_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08138__S _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14480_/A sky130_fd_sc_hd__buf_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11673_ _11673_/A _11758_/C vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__xnor2_1
XFILLER_169_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14664__A _14681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13412_ _13401_/A _13747_/B _13411_/X vssd1 vssd1 vccd1 vccd1 _13448_/A sky130_fd_sc_hd__a21bo_1
XANTENNA_input90_A x_i_5[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ _10622_/A _10622_/B _10623_/X vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__a21oi_1
XFILLER_139_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14392_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14392_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12963__A1 _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11800__B _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ _13373_/A _13343_/B vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__xor2_4
XFILLER_182_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10555_ _15262_/Q _15295_/Q vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__or2b_1
XFILLER_155_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13274_ _13274_/A _13274_/B _13274_/C vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__and3_1
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10486_ _10486_/A _10486_/B vssd1 vssd1 vccd1 vccd1 _14904_/D sky130_fd_sc_hd__xnor2_1
X_15013_ _15435_/CLK _15013_/D _14049_/Y vssd1 vssd1 vccd1 vccd1 _15013_/Q sky130_fd_sc_hd__dfrtp_1
X_12225_ _12219_/A _12219_/B _12222_/X _12224_/X vssd1 vssd1 vccd1 vccd1 _12268_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12156_ _12156_/A _12156_/B _12556_/B vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__and3_1
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output344_A output344/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11107_ _11107_/A _11107_/B vssd1 vssd1 vccd1 vccd1 _11107_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_190_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12087_ _12087_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nor2_1
Xrepeater907 repeater908/X vssd1 vssd1 vccd1 vccd1 _07738_/A1 sky130_fd_sc_hd__buf_4
Xrepeater918 input190/X vssd1 vssd1 vccd1 vccd1 _07695_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater929 input176/X vssd1 vssd1 vccd1 vccd1 _07822_/A1 sky130_fd_sc_hd__clkbuf_2
X_11038_ _14926_/Q _14992_/Q vssd1 vssd1 vccd1 vccd1 _11039_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output511_A output511/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__B _15310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14839__A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater661_A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15777_ _15777_/CLK _15777_/D _14856_/Y vssd1 vssd1 vccd1 vccd1 _15777_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12989_ _13688_/A _13688_/B _12976_/C _12988_/X _12912_/B vssd1 vssd1 vccd1 vccd1
+ _12989_/X sky130_fd_sc_hd__o311a_1
XANTENNA_repeater759_A _15643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14728_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14659_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater926_A repeater927/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14574__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08180_ _11707_/A _11617_/A vssd1 vssd1 vccd1 vccd1 _08185_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08572__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12954__A1 _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13918__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12822__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput267 _11104_/Y vssd1 vssd1 vccd1 vccd1 y_i_0[16] sky130_fd_sc_hd__buf_2
XFILLER_88_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput278 output278/A vssd1 vssd1 vccd1 vccd1 y_i_1[10] sky130_fd_sc_hd__buf_2
XFILLER_47_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput289 _15648_/Q vssd1 vssd1 vccd1 vccd1 y_i_1[5] sky130_fd_sc_hd__buf_2
XFILLER_88_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11438__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ _15709_/Q _14987_/Q vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__or2_1
XFILLER_4_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09703_ _09824_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _15713_/D sky130_fd_sc_hd__xnor2_1
XFILLER_68_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07895_ _07895_/A vssd1 vssd1 vccd1 vccd1 _15320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14749__A _14750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09634_ _15563_/Q vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11693__A1 _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ _15434_/Q _15418_/Q vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07649__A0 _15441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08516_ _08516_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _08681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09496_ _15526_/Q _15510_/Q vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__and2_1
XFILLER_54_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ _13203_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_759 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14484__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__A _15438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08378_ _12921_/A _12810_/A vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_762 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ _15128_/Q _15161_/Q _10336_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _15082_/Q _15247_/Q vssd1 vssd1 vccd1 vccd1 _10273_/A sky130_fd_sc_hd__or2b_1
X_12010_ _12011_/A _12011_/B _12009_/Y vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__o21bai_1
XFILLER_151_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12451__B _12451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input242_A x_r_6[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13961_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13961_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14659__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07888__A0 _15323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12912_/A _12912_/B vssd1 vssd1 vccd1 vccd1 _13677_/C sky130_fd_sc_hd__nand2_4
XFILLER_47_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15700_ _15700_/CLK _15700_/D _14775_/Y vssd1 vssd1 vccd1 vccd1 _15700_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_111_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13892_ _15340_/Q _15324_/Q _13891_/X vssd1 vssd1 vccd1 vccd1 _13893_/B sky130_fd_sc_hd__a21oi_1
XFILLER_206_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15631_ _15680_/CLK _15631_/D _14703_/Y vssd1 vssd1 vccd1 vccd1 _15631_/Q sky130_fd_sc_hd__dfrtp_1
X_12843_ _12843_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _12845_/A sky130_fd_sc_hd__nand2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _15563_/CLK _15562_/D _14629_/Y vssd1 vssd1 vccd1 vccd1 _15562_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A _12774_/B vssd1 vssd1 vccd1 vccd1 _15628_/D sky130_fd_sc_hd__xnor2_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14513_/Y sky130_fd_sc_hd__inv_2
X_11725_ _15730_/Q _11725_/B vssd1 vssd1 vccd1 vccd1 _11725_/X sky130_fd_sc_hd__and2_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ _15493_/CLK _15493_/D _14556_/Y vssd1 vssd1 vccd1 vccd1 _15493_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14394__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14444_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11656_ _11654_/A _12533_/A _11655_/X vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__a21o_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07500__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output294_A output294/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10607_ _15260_/Q _15293_/Q _10606_/B vssd1 vssd1 vccd1 vccd1 _10609_/C sky130_fd_sc_hd__a21o_1
X_14375_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14375_/Y sky130_fd_sc_hd__inv_2
X_11587_ _11898_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13326_ _14920_/Q _13327_/B vssd1 vssd1 vccd1 vccd1 _13380_/A sky130_fd_sc_hd__and2_1
XFILLER_183_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10538_ _10538_/A _10543_/A vssd1 vssd1 vccd1 vccd1 _15028_/D sky130_fd_sc_hd__nor2_1
XANTENNA_output461_A output461/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13257_ _13257_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _13258_/B sky130_fd_sc_hd__and2_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10469_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__and3_1
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12208_ _12208_/A _12207_/Y vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__or2b_1
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _13189_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13263_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ _12139_/A _12187_/A vssd1 vssd1 vccd1 vccd1 _12141_/C sky130_fd_sc_hd__xnor2_1
XFILLER_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater704 _07644_/S vssd1 vssd1 vccd1 vccd1 _07632_/S sky130_fd_sc_hd__buf_8
XFILLER_29_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater715 _15704_/Q vssd1 vssd1 vccd1 vccd1 output382/A sky130_fd_sc_hd__buf_4
XFILLER_38_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater726 _15690_/Q vssd1 vssd1 vccd1 vccd1 output350/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater737 _15665_/Q vssd1 vssd1 vccd1 vccd1 output323/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater748 _15654_/Q vssd1 vssd1 vccd1 vccd1 repeater748/X sky130_fd_sc_hd__buf_2
XANTENNA__14569__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater759 _15643_/Q vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ _07680_/A vssd1 vssd1 vccd1 vccd1 _15426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09350_ _15397_/Q _09351_/B _09351_/C vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__a21o_1
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08301_ _08293_/Y _11545_/A _08291_/Y _08292_/Y _08300_/Y vssd1 vssd1 vccd1 vccd1
+ _08301_/X sky130_fd_sc_hd__a221o_1
X_09281_ _15399_/Q _15383_/Q vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__and2_1
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08843__A2 _15331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07410__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__B _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ _11469_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10337__A _15129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__B_N _08968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07803__A0 _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08094_ _08094_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08120_/C sky130_fd_sc_hd__xor2_2
XFILLER_109_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07646__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1063 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08996_ _15368_/Q _15352_/Q vssd1 vssd1 vccd1 vccd1 _08996_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07947_ _15251_/Q _15284_/Q vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__or2_1
XANTENNA__14479__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07878_ _15328_/Q _07878_/A1 _07892_/S vssd1 vssd1 vccd1 vccd1 _07879_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07381__A _07434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _09617_/A _09617_/B vssd1 vssd1 vccd1 vccd1 _15182_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_838 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ _15432_/Q _15416_/Q vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__xnor2_2
XFILLER_203_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1064 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__B1 _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ _09479_/A _09484_/A vssd1 vssd1 vccd1 vccd1 _09529_/A sky130_fd_sc_hd__or2_1
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11631__A _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _11510_/A _11456_/A vssd1 vssd1 vccd1 vccd1 _11537_/A sky130_fd_sc_hd__or2b_1
XFILLER_180_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ _12490_/A vssd1 vssd1 vccd1 vccd1 _15655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ _11876_/A _11977_/A vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__xor2_2
XANTENNA_input192_A x_r_3[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14160_/Y sky130_fd_sc_hd__inv_2
X_11372_ _11372_/A _11372_/B _11372_/C vssd1 vssd1 vccd1 vccd1 _11375_/B sky130_fd_sc_hd__and3_1
XFILLER_124_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_946 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13111_ _13153_/A _12859_/C _13319_/A vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__mux2_1
X_10323_ _15126_/Q _15159_/Q vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__nand2_1
X_14091_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14091_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input53_A x_i_3[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _13042_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _13042_/X sky130_fd_sc_hd__or2_1
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10254_ _10253_/A _10253_/B _11411_/B vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__a21o_1
XFILLER_191_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ _10183_/A _10854_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _10187_/A sky130_fd_sc_hd__o21ai_1
XFILLER_121_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14389__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14993_ _15027_/CLK _14993_/D _14027_/Y vssd1 vssd1 vccd1 vccd1 _14993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11806__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13944_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13944_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _15334_/Q _15318_/Q vssd1 vssd1 vccd1 vccd1 _13875_/X sky130_fd_sc_hd__and2_1
XFILLER_19_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output307_A output307/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15614_ _15689_/CLK _15614_/D _14685_/Y vssd1 vssd1 vccd1 vccd1 _15614_/Q sky130_fd_sc_hd__dfrtp_2
X_12826_ _12826_/A _12826_/B vssd1 vssd1 vccd1 vccd1 _12882_/A sky130_fd_sc_hd__xnor2_1
XFILLER_201_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15545_ _15568_/CLK _15545_/D _14611_/Y vssd1 vssd1 vccd1 vccd1 _15545_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12779_/A _12779_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__xor2_2
XFILLER_188_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12637__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_135_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15525_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11708_ _11709_/A _11709_/B _11709_/C vssd1 vssd1 vccd1 vccd1 _11710_/A sky130_fd_sc_hd__a21oi_1
XFILLER_203_696 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15476_ _15511_/CLK _15476_/D _14538_/Y vssd1 vssd1 vccd1 vccd1 _15476_/Q sky130_fd_sc_hd__dfrtp_4
X_12688_ _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _12690_/C sky130_fd_sc_hd__xnor2_1
XFILLER_175_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14427_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11639_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__xor2_1
XANTENNA_repeater624_A _11111_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14852__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13309_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14289_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14289_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_532 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08850_ _08855_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08936_/B sky130_fd_sc_hd__or2_1
XFILLER_123_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07801_ _15366_/Q _07801_/A1 _07803_/S vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _13883_/A _08778_/B _08780_/X vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14299__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater534 _13706_/X vssd1 vssd1 vccd1 vccd1 _15699_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater545 _10806_/Y vssd1 vssd1 vccd1 vccd1 output403/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11716__A _11728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _15400_/Q _07732_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater556 _11289_/Y vssd1 vssd1 vccd1 vccd1 repeater556/X sky130_fd_sc_hd__buf_4
XFILLER_66_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater567 _10789_/X vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__buf_2
Xrepeater578 repeater579/X vssd1 vssd1 vccd1 vccd1 output431/A sky130_fd_sc_hd__buf_4
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater589 _10769_/Y vssd1 vssd1 vccd1 vccd1 output397/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08728__C _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _15434_/Q _07663_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09402_ _09401_/Y _15395_/Q _09400_/B vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13931__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07594_ _15468_/Q input80/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09333_ _15409_/Q _15393_/Q vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__and2_1
XFILLER_52_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_126_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15500_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_392 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _15506_/Q _15490_/Q vssd1 vssd1 vccd1 vccd1 _09266_/A sky130_fd_sc_hd__or2b_1
XFILLER_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12266__B _12564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08215_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09195_ _09195_/A _09667_/A vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__nand2_1
XFILLER_194_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _15017_/Q vssd1 vssd1 vccd1 vccd1 _12254_/A sky130_fd_sc_hd__buf_4
XFILLER_153_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ _12055_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09575__B _15420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14912__D _14912_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13876__A2 _15317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ _15366_/Q _15350_/Q vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__and2b_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ _11990_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14002__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12300__A2 _12564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10941_ _10941_/A vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08000__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13660_ _13816_/A _13816_/B vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__xnor2_4
X_10872_ _10872_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _11109_/A sky130_fd_sc_hd__nand2_2
XANTENNA_input205_A x_r_4[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12611_ _12496_/A _12496_/B _12610_/B vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__a21oi_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15764_/CLK sky130_fd_sc_hd__clkbuf_16
X_13591_ _13591_/A _13591_/B vssd1 vssd1 vccd1 vccd1 _15087_/D sky130_fd_sc_hd__xnor2_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15341_/CLK _15330_/D _14384_/Y vssd1 vssd1 vccd1 vccd1 _15330_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12536_/A _12537_/A _12536_/B _12538_/X _11788_/B vssd1 vssd1 vccd1 vccd1
+ _12543_/B sky130_fd_sc_hd__a311o_1
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15261_ _15268_/CLK _15261_/D _14311_/Y vssd1 vssd1 vccd1 vccd1 _15261_/Q sky130_fd_sc_hd__dfrtp_1
X_12473_ _12460_/Y _12465_/B _12461_/A vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__a21o_1
XFILLER_177_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14672__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14212_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14212_/Y sky130_fd_sc_hd__inv_2
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _15740_/D sky130_fd_sc_hd__xor2_2
XFILLER_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _15192_/CLK _15192_/D _14237_/Y vssd1 vssd1 vccd1 vccd1 _15192_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14143_/Y sky130_fd_sc_hd__inv_2
X_11355_ _11355_/A _11355_/B vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_180_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _10443_/A _10306_/B vssd1 vssd1 vccd1 vccd1 _15778_/D sky130_fd_sc_hd__xnor2_2
XFILLER_113_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14074_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11286_ _11286_/A vssd1 vssd1 vccd1 vccd1 _11286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13025_ _13025_/A _13025_/B vssd1 vssd1 vccd1 vccd1 _13036_/A sky130_fd_sc_hd__nor2_1
X_10237_ _10235_/Y _10237_/B vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__and2b_1
XFILLER_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _10168_/A _10168_/B _10850_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__and3_1
XFILLER_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output424_A output424/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _15301_/Q _15136_/Q vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__or2b_1
X_14976_ _15249_/CLK _14976_/D _14009_/Y vssd1 vssd1 vccd1 vccd1 _14976_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13927_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13927_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater574_A _11377_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14847__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13858_ _13858_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13859_/A sky130_fd_sc_hd__nor2_1
XFILLER_179_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater741_A _15659_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _13677_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_108_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15774_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_repeater839_A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _13789_/A _13863_/A vssd1 vssd1 vccd1 vccd1 _15706_/D sky130_fd_sc_hd__xor2_1
XFILLER_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15528_ _15528_/CLK _15528_/D _14593_/Y vssd1 vssd1 vccd1 vccd1 _15528_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15459_ _15700_/CLK _15459_/D _14520_/Y vssd1 vssd1 vccd1 vccd1 _15459_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14582__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08000_ _11876_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _08009_/C sky130_fd_sc_hd__xor2_2
XFILLER_50_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08982__A1 _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _15231_/Q _15198_/Q vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__or2b_1
XFILLER_171_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ _08900_/X _08907_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13926__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09882_ _15187_/Q _09881_/Y _09877_/B vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__a21o_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07924__A _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08832_/A _08832_/B _13908_/A vssd1 vssd1 vccd1 vccd1 _08836_/B sky130_fd_sc_hd__a21oi_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11446__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08764_ _08766_/B _08764_/B vssd1 vssd1 vccd1 vccd1 _15070_/D sky130_fd_sc_hd__nor2_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07715_ _07715_/A vssd1 vssd1 vccd1 vccd1 _15409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08695_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__xor2_2
XFILLER_199_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14757__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07695_/S sky130_fd_sc_hd__buf_8
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07577_ _15476_/Q input73/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07578_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09316_ _09377_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _15128_/D sky130_fd_sc_hd__xor2_2
XANTENNA__12708__C _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_896 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ _09247_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__and2_1
XANTENNA__07473__A1 _07473_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14492__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09586__A _15438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09178_ _09652_/A _09178_/B vssd1 vssd1 vccd1 vccd1 _15292_/D sky130_fd_sc_hd__xnor2_1
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15738__D _15738_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08129_ _11832_/A _11687_/A vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__xor2_2
XFILLER_31_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ _11140_/A _11140_/B vssd1 vssd1 vccd1 vccd1 _11140_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_107_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11071_ _11072_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11071_/X sky130_fd_sc_hd__xor2_1
XANTENNA_input155_A x_r_1[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput101 x_i_6[11] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 x_i_6[7] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_2
X_10022_ _15204_/Q _15105_/Q vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput123 x_i_7[2] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput134 x_r_0[12] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_2
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 x_r_0[8] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__clkbuf_2
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput156 x_r_1[3] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_2
Xinput167 x_r_2[13] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_2
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14830_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14830_/Y sky130_fd_sc_hd__inv_2
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 x_r_2[9] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput189 x_r_3[4] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A x_i_0[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11973_ _12031_/A _12031_/B vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__xnor2_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14761_/Y sky130_fd_sc_hd__inv_2
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14667__A _14681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _10924_/A _10924_/B _11124_/B vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__and3_1
X_13712_ _13712_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14692_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08665__A _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11803__B _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _10854_/A _10854_/B _10182_/B vssd1 vssd1 vccd1 vccd1 _10856_/B sky130_fd_sc_hd__a21oi_1
X_13643_ _08757_/A _13809_/B _13642_/X vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__a21oi_2
XFILLER_73_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08384__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _13574_/A _13574_/B vssd1 vssd1 vccd1 vccd1 _15605_/D sky130_fd_sc_hd__xor2_2
XFILLER_73_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ _10786_/A _10786_/B vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__nor2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12525_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__xor2_1
XFILLER_160_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15313_ _15569_/CLK _15313_/D _14366_/Y vssd1 vssd1 vccd1 vccd1 _15313_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12456_ _12456_/A _12456_/B _12456_/C _12456_/D vssd1 vssd1 vccd1 vccd1 _12458_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15244_ _15764_/CLK _15244_/D _14293_/Y vssd1 vssd1 vccd1 vccd1 _15244_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output374_A output374/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _10235_/Y _11406_/B _10237_/B vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__o21ai_2
X_15175_ _15175_/CLK _15175_/D _14220_/Y vssd1 vssd1 vccd1 vccd1 _15175_/Q sky130_fd_sc_hd__dfrtp_1
X_12387_ _12586_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__and2b_1
XFILLER_158_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12633__B_N _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _11338_/A vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14057_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14057_/Y sky130_fd_sc_hd__inv_2
X_11269_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11269_/Y sky130_fd_sc_hd__nor2_2
XFILLER_122_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _13008_/A _13008_/B _13008_/C vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__and3_1
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater691_A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater789_A _15603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ _15809_/CLK _14959_/D _13991_/Y vssd1 vssd1 vccd1 vccd1 _14959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater956_A input140/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14577__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _15514_/Q input30/X _07536_/S vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08480_ _14915_/Q vssd1 vssd1 vccd1 vccd1 _13381_/B sky130_fd_sc_hd__buf_6
XFILLER_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07431_ _07431_/A vssd1 vssd1 vccd1 vccd1 _15548_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09101_ _15501_/Q _15485_/Q vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__xnor2_2
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07455__A1 _07455_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09032_ _09031_/A _09031_/B _13614_/B vssd1 vssd1 vccd1 vccd1 _09038_/B sky130_fd_sc_hd__a21o_1
XFILLER_191_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _09932_/X _09939_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A x_i_0[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _15758_/D sky130_fd_sc_hd__xnor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08816_ _15344_/Q _15328_/Q vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__or2b_1
X_09796_ _09795_/A _09795_/C _09795_/B vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__o21a_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ _08707_/Y _08712_/Y _08744_/X _08746_/X vssd1 vssd1 vccd1 vccd1 _08750_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_90_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14487__A _14488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_944 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08678_ _12780_/A _08478_/A _08677_/Y vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__a21oi_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08485__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__B _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ _07629_/A vssd1 vssd1 vccd1 vccd1 _15451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ _15270_/Q _15171_/Q vssd1 vssd1 vccd1 vccd1 _10642_/A sky130_fd_sc_hd__or2_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _10571_/A _10577_/A vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12735__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12310_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13290_ _13290_/A _13700_/A vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__and2_1
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12241_ _12239_/Y _12241_/B vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__and2b_1
XFILLER_154_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _12171_/B _12172_/B vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__and2b_1
XFILLER_135_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _11124_/A _11124_/C _11124_/B vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_43_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11054_ _11052_/Y _11054_/B vssd1 vssd1 vccd1 vccd1 _11327_/A sky130_fd_sc_hd__and2b_1
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_693 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ _10003_/A _10003_/B _10004_/X vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__a21oi_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14813_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_922 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15793_ _15795_/CLK _15793_/D _14873_/Y vssd1 vssd1 vccd1 vccd1 _15793_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14397__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_101_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14744_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ _12308_/S _12228_/A vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__xor2_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08395__A _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08331__C1 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07685__A1 input180/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ _14962_/Q _14896_/Q vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11887_ _11887_/A _11887_/B vssd1 vssd1 vccd1 vccd1 _11954_/A sky130_fd_sc_hd__xnor2_1
X_14675_ _14675_/A vssd1 vssd1 vccd1 vccd1 _14675_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10838_ _15309_/Q _15144_/Q vssd1 vssd1 vccd1 vccd1 _10839_/C sky130_fd_sc_hd__or2b_1
X_13626_ _15378_/Q _15362_/Q vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__and2_1
XFILLER_38_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output491_A _15613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09582__A_N _15437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_116_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__A1 _07437_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10769_ _11283_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10769_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_125_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13557_ _15766_/Q _13563_/B vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12508_ _12508_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__and2_1
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13488_ _13505_/A _13505_/B vssd1 vssd1 vccd1 vccd1 _13790_/A sky130_fd_sc_hd__xor2_2
XFILLER_195_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ _12427_/B _12439_/B vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__and2b_1
X_15227_ _15501_/CLK _15227_/D _14275_/Y vssd1 vssd1 vccd1 vccd1 _15227_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater704_A _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14860__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput405 output405/A vssd1 vssd1 vccd1 vccd1 y_r_0[2] sky130_fd_sc_hd__buf_2
XFILLER_172_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput416 _15589_/Q vssd1 vssd1 vccd1 vccd1 y_r_1[12] sky130_fd_sc_hd__buf_2
Xoutput427 output427/A vssd1 vssd1 vccd1 vccd1 y_r_1[7] sky130_fd_sc_hd__buf_2
X_15158_ _15434_/CLK _15158_/D _14202_/Y vssd1 vssd1 vccd1 vccd1 _15158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput438 output438/A vssd1 vssd1 vccd1 vccd1 y_r_2[1] sky130_fd_sc_hd__buf_2
Xoutput449 _15605_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[11] sky130_fd_sc_hd__buf_2
XFILLER_153_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14109_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07980_ _15796_/Q vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15089_ _15712_/CLK _15089_/D _14129_/Y vssd1 vssd1 vccd1 vccd1 _15089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ _09648_/A _09648_/B _09649_/X vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ _08715_/B _08715_/A vssd1 vssd1 vccd1 vccd1 _08601_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _09581_/A vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08532_ _14913_/Q vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__buf_4
XFILLER_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14100__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08463_ _08451_/A _08451_/B _08466_/A vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__a21o_1
XFILLER_35_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ _15556_/Q input57/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08394_ _12654_/A _08396_/C vssd1 vssd1 vccd1 vccd1 _08434_/B sky130_fd_sc_hd__nand2_1
XFILLER_189_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07428__A1 _07428_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15576_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09013_/Y _09015_/B vssd1 vssd1 vccd1 vccd1 _13610_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__14770__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14920__D _14920_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07600__A1 _07600_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12290__A _12291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09917_ _15225_/Q _15192_/Q vssd1 vssd1 vccd1 vccd1 _09918_/C sky130_fd_sc_hd__or2b_1
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_97_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _09848_/A _09848_/B _09848_/C vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__and3_1
XFILLER_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _15432_/Q _15416_/Q _09778_/B vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11878_/A _11877_/A vssd1 vssd1 vccd1 vccd1 _11811_/B sky130_fd_sc_hd__xor2_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A _12859_/C vssd1 vssd1 vccd1 vccd1 _12791_/C sky130_fd_sc_hd__xnor2_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A x_i_7[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14010__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11842_/C _11849_/B _11928_/A vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07667__A1 input252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11758_/C sky130_fd_sc_hd__xor2_1
X_14460_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14460_/Y sky130_fd_sc_hd__inv_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13411_ _13411_/A _13399_/A vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__or2b_1
X_10623_ _15265_/Q _15298_/Q vssd1 vssd1 vccd1 vccd1 _10623_/X sky130_fd_sc_hd__and2_1
XFILLER_186_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14391_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14391_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15220_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13342_ _13247_/A _13247_/B _13245_/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13343_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_210_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input83_A x_i_5[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10554_ _10554_/A vssd1 vssd1 vccd1 vccd1 _15030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_944 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _13273_/A _13273_/B vssd1 vssd1 vccd1 vccd1 _13274_/C sky130_fd_sc_hd__xnor2_1
XFILLER_185_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10485_ _10484_/A _10484_/B _10374_/B vssd1 vssd1 vccd1 vccd1 _10486_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14680__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15012_ _15663_/CLK _15012_/D _14048_/Y vssd1 vssd1 vccd1 vccd1 _15012_/Q sky130_fd_sc_hd__dfrtp_1
X_12224_ _12156_/B _12223_/X _12560_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12224_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12155_ _12220_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__or2_2
XFILLER_118_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _14955_/Q _15809_/Q _10860_/Y _10861_/Y vssd1 vssd1 vccd1 vccd1 _11107_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12086_ _12086_/A _12086_/B _12086_/C vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__and3_1
XFILLER_111_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output337_A _11305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15107_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater908 input211/X vssd1 vssd1 vccd1 vccd1 repeater908/X sky130_fd_sc_hd__buf_2
Xrepeater919 input19/X vssd1 vssd1 vccd1 vccd1 _07510_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11037_ _14926_/Q _14992_/Q vssd1 vssd1 vccd1 vccd1 _11039_/A sky130_fd_sc_hd__or2_1
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12884__D1 _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output504_A output504/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15661__D _15661_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15776_ _15777_/CLK _15776_/D _14855_/Y vssd1 vssd1 vccd1 vccd1 _15776_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12910_/A _12985_/B _12910_/C _12986_/B _13677_/A vssd1 vssd1 vccd1 vccd1
+ _12988_/X sky130_fd_sc_hd__a32o_1
XFILLER_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09014__A _15373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14727_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14727_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11939_ _11783_/A _11783_/B _11793_/X _11794_/X _12406_/A vssd1 vssd1 vccd1 vccd1
+ _11940_/B sky130_fd_sc_hd__o311a_1
XFILLER_178_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater654_A _07957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14855__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14658_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13609_ _15372_/Q _15356_/Q _13608_/X vssd1 vssd1 vccd1 vccd1 _13610_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater821_A input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14589_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14589_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08572__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15561_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12954__A2 _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_988 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07830__A1 _07830_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14590__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12822__B _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11719__A _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput268 _11020_/Y vssd1 vssd1 vccd1 vccd1 y_i_0[1] sky130_fd_sc_hd__buf_2
XANTENNA__07916__B _15509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput279 output279/A vssd1 vssd1 vccd1 vccd1 y_i_1[11] sky130_fd_sc_hd__buf_2
XFILLER_88_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07594__A0 _15468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07408__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _15709_/Q _14987_/Q vssd1 vssd1 vccd1 vccd1 _11353_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_79_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 _15724_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13934__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ _09696_/A _09698_/B _09696_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__a21boi_1
XFILLER_114_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07894_ _15320_/Q _07894_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07895_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09633_ _09633_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _15302_/D sky130_fd_sc_hd__nor2_1
XANTENNA__11693__A2 _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09564_ _09562_/Y _09564_/B vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__nand2b_1
XFILLER_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ _13046_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07649__A1 input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _09495_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _15252_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__14765__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08763__A _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ _15048_/Q vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__buf_4
XANTENNA__14915__D _14915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09594__A _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10270_ _10270_/A vssd1 vssd1 vccd1 vccd1 _15770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15746__D _15746_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14005__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08845__A_N _15348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__B _11348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input235_A x_r_6[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_803 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13960_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12330__A0 _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12911_ _12985_/B _12910_/C _12910_/A vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07888__A1 _07888_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13563__B _13563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13891_ _15340_/Q _15324_/Q _13890_/B vssd1 vssd1 vccd1 vccd1 _13891_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15630_ _15680_/CLK _15630_/D _14701_/Y vssd1 vssd1 vccd1 vccd1 _15630_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12842_ _15761_/Q _13539_/B vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__xnor2_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/CLK _15561_/D _14628_/Y vssd1 vssd1 vccd1 vccd1 _15561_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_203_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12894__S _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12843_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _12774_/B sky130_fd_sc_hd__xnor2_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14675__A _14675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14512_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11724_ _12537_/A vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15572_/CLK _15492_/D _14555_/Y vssd1 vssd1 vccd1 vccd1 _15492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11655_ _12534_/B _15729_/Q vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__and2b_1
X_14443_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14443_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _14996_/D sky130_fd_sc_hd__xnor2_1
XFILLER_196_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11586_ _11530_/A _11530_/B _11585_/X vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__a21oi_1
XFILLER_167_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14374_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14374_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output287_A output287/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _13325_/A _13325_/B vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__xor2_1
X_10537_ _10536_/A _10536_/C _10604_/A vssd1 vssd1 vccd1 vccd1 _10543_/A sky130_fd_sc_hd__a21oi_1
XFILLER_156_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_796 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10468_ _15161_/Q _15128_/Q vssd1 vssd1 vccd1 vccd1 _10469_/C sky130_fd_sc_hd__or2b_1
X_13256_ _13257_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__nor2_1
X_12207_ _12207_/A _12207_/B _12207_/C vssd1 vssd1 vccd1 vccd1 _12207_/Y sky130_fd_sc_hd__nand3_1
X_13187_ _13187_/A _13187_/B vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__xnor2_1
X_10399_ _15107_/Q _15206_/Q vssd1 vssd1 vccd1 vccd1 _10400_/C sky130_fd_sc_hd__or2b_1
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _12074_/A _12074_/B _12073_/A vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09009__A _15372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater705 _07575_/S vssd1 vssd1 vccd1 vccd1 _07589_/S sky130_fd_sc_hd__buf_4
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12069_ _12071_/A _12144_/A _12247_/A _11987_/X _12254_/A vssd1 vssd1 vccd1 vccd1
+ _12073_/A sky130_fd_sc_hd__o2111a_1
Xrepeater716 _15703_/Q vssd1 vssd1 vccd1 vccd1 output381/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater727 _15685_/Q vssd1 vssd1 vccd1 vccd1 output361/A sky130_fd_sc_hd__clkbuf_2
Xrepeater738 _15663_/Q vssd1 vssd1 vccd1 vccd1 output321/A sky130_fd_sc_hd__clkbuf_2
Xrepeater749 _15653_/Q vssd1 vssd1 vccd1 vccd1 output278/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07752__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater771_A repeater772/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09000__A_N _15369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15759_ _15761_/CLK _15759_/D _14837_/Y vssd1 vssd1 vccd1 vccd1 _15759_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14585__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ _11678_/A _11707_/A _11687_/A _11658_/A _08299_/X vssd1 vssd1 vccd1 vccd1
+ _08300_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_178_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07898__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _15398_/Q _09275_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07500__A0 _15514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08231_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__xnor2_1
XFILLER_193_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08093_ _08101_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13929__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07803__A1 input227/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08995_ _08993_/Y _08995_/B vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__nand2b_1
XFILLER_134_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07946_ _15251_/Q _15284_/Q vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08758__A _15317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _07877_/A vssd1 vssd1 vccd1 vccd1 _15329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _09615_/A _09615_/B _09809_/A vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__o21a_1
XFILLER_18_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09547_ _09547_/A _09547_/B vssd1 vssd1 vccd1 vccd1 _15170_/D sky130_fd_sc_hd__nor2_1
XANTENNA__14495__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08493__A _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09478_ _15538_/Q _15522_/Q vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__and2b_1
XFILLER_93_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ _08429_/A _08429_/B _08427_/Y vssd1 vssd1 vccd1 vccd1 _08430_/B sky130_fd_sc_hd__or3b_1
XFILLER_180_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09643__A_N _15566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11440_ _11898_/A _11797_/A vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09101__B _15485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_780 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11371_ _11372_/A _11372_/C _11372_/B vssd1 vssd1 vccd1 vccd1 _11373_/A sky130_fd_sc_hd__a21oi_1
XFILLER_152_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input185_A x_r_3[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12743__A _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10322_ _15126_/Q _15159_/Q vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__or2_1
XFILLER_3_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13110_ _13381_/B vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__inv_2
XFILLER_152_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14090_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13558__B _13558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13041_ _13041_/A _13041_/B vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10253_ _10253_/A _10253_/B _11411_/B vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__and3_1
XFILLER_65_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A x_i_2[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _15150_/Q _15315_/Q vssd1 vssd1 vccd1 vccd1 _10184_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09023__A_N _15373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14992_ _15027_/CLK _14992_/D _14026_/Y vssd1 vssd1 vccd1 vccd1 _14992_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11806__B _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13943_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13943_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11511__D1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ _13874_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _15054_/D sky130_fd_sc_hd__xnor2_1
XFILLER_189_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15613_ _15649_/CLK _15613_/D _14684_/Y vssd1 vssd1 vccd1 vccd1 _15613_/Q sky130_fd_sc_hd__dfrtp_1
X_12825_ _12825_/A _12825_/B vssd1 vssd1 vccd1 vccd1 _12826_/B sky130_fd_sc_hd__xnor2_1
XFILLER_203_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15563_/CLK _15544_/D _14610_/Y vssd1 vssd1 vccd1 vccd1 _15544_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_163_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12683_/A _12754_/Y _12755_/Y vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__o21ai_2
XFILLER_199_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A _11707_/B vssd1 vssd1 vccd1 vccd1 _11709_/C sky130_fd_sc_hd__xnor2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15475_ _15509_/CLK _15475_/D _14537_/Y vssd1 vssd1 vccd1 vccd1 _15475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ _12687_/A _12759_/A vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__xnor2_2
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14426_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14426_/Y sky130_fd_sc_hd__inv_2
X_11638_ _11638_/A _11638_/B vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14357_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14357_/Y sky130_fd_sc_hd__inv_2
X_11569_ _11569_/A _11569_/B _11569_/C vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__and3_1
XANTENNA_repeater617_A _11169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__A0 _15368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__or3_1
XFILLER_144_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14288_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14288_/Y sky130_fd_sc_hd__inv_2
X_13239_ _13333_/B _13239_/B vssd1 vssd1 vccd1 vccd1 _13240_/C sky130_fd_sc_hd__or2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater986_A input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _07800_/A vssd1 vssd1 vccd1 vccd1 _15367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08780_ _15337_/Q _15321_/Q vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__and2b_1
XFILLER_211_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A vssd1 vssd1 vccd1 vccd1 _15401_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater535 _13826_/Y vssd1 vssd1 vccd1 vccd1 _15666_/D sky130_fd_sc_hd__clkbuf_2
Xrepeater546 _12575_/X vssd1 vssd1 vccd1 vccd1 _15677_/D sky130_fd_sc_hd__buf_4
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater557 _11218_/X vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10620__B _15297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater568 _11379_/X vssd1 vssd1 vccd1 vccd1 output433/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater579 _11373_/Y vssd1 vssd1 vccd1 vccd1 repeater579/X sky130_fd_sc_hd__buf_2
X_07662_ _07662_/A vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08728__D _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09401_ _15411_/Q vssd1 vssd1 vccd1 vccd1 _09401_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07593_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07644_/S sky130_fd_sc_hd__buf_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _09332_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _15131_/D sky130_fd_sc_hd__xor2_4
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _09265_/A _09265_/B vssd1 vssd1 vccd1 vccd1 _15247_/D sky130_fd_sc_hd__xor2_1
XFILLER_179_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08214_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__xor2_1
XFILLER_166_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09226__B1 _09224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09194_ _15572_/Q _15552_/Q vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__or2b_1
XFILLER_53_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08145_ _12204_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09777__A1 _15431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08076_ _11806_/C _08094_/A _08076_/C vssd1 vssd1 vccd1 vccd1 _08090_/A sky130_fd_sc_hd__or3_1
XFILLER_174_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09872__A _15187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08978_ _15349_/Q vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__inv_2
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07929_ _15185_/Q _15218_/Q vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _10938_/X _10945_/B vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__and2b_1
XFILLER_57_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08000__B _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10871_ _14957_/Q _14891_/Q vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12738__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12610_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _15689_/D sky130_fd_sc_hd__xnor2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input100_A x_i_6[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _15610_/D sky130_fd_sc_hd__xnor2_1
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _15731_/Q _12541_/B vssd1 vssd1 vccd1 vccd1 _12543_/A sky130_fd_sc_hd__or2_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15260_ _15561_/CLK _15260_/D _14310_/Y vssd1 vssd1 vccd1 vccd1 _15260_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_196_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12472_ _12472_/A vssd1 vssd1 vccd1 vccd1 _12604_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14211_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11423_ _11421_/A _11421_/B _11422_/X vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__a21o_1
X_15191_ _15192_/CLK _15191_/D _14236_/Y vssd1 vssd1 vccd1 vccd1 _15191_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07779__A0 _15377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11354_ _15743_/Q _15021_/Q _11147_/Y _11248_/A vssd1 vssd1 vccd1 vccd1 _11355_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14142_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10305_ _10301_/A _10298_/Y _10300_/B vssd1 vssd1 vccd1 vccd1 _10306_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__08991__A2 _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11285_ _11283_/X _11287_/C vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__and2b_2
X_14073_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14073_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _13023_/B _13023_/C _13023_/A vssd1 vssd1 vccd1 vccd1 _13100_/B sky130_fd_sc_hd__a21o_1
X_10236_ _15077_/Q _15242_/Q vssd1 vssd1 vccd1 vccd1 _10237_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10167_ _10167_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__nor2_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08398__A _15045_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14975_ _15249_/CLK _14975_/D _14008_/Y vssd1 vssd1 vccd1 vccd1 _14975_/Q sky130_fd_sc_hd__dfrtp_1
X_10098_ _10098_/A _10434_/A vssd1 vssd1 vccd1 vccd1 _14986_/D sky130_fd_sc_hd__xnor2_1
XFILLER_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output417_A output417/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13926_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13926_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13857_ _14982_/Q vssd1 vssd1 vccd1 vccd1 _13858_/A sky130_fd_sc_hd__inv_2
XFILLER_63_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08845__B _15332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _13057_/A _13056_/C _13057_/B _12807_/Y vssd1 vssd1 vccd1 vccd1 _12809_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13788_ _13788_/A _13788_/B vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _15527_/CLK _15527_/D _14592_/Y vssd1 vssd1 vccd1 vccd1 _15527_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12739_ _12970_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14863__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater734_A _15672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15458_ _15472_/CLK _15458_/D _14519_/Y vssd1 vssd1 vccd1 vccd1 _15458_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14409_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater901_A repeater902/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15389_ _15411_/CLK _15389_/D _14447_/Y vssd1 vssd1 vccd1 vccd1 _15389_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09950_ _15198_/Q _15231_/Q vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1020 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08901_ _08900_/A _08900_/B _08959_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _15220_/Q vssd1 vssd1 vccd1 vccd1 _09881_/Y sky130_fd_sc_hd__inv_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08832_ _08832_/A _08832_/B _13908_/A vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__and3_1
XFILLER_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07924__B _15541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14103__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07416__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_942 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08763_ _15333_/Q _08763_/B _13874_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__and3_1
XFILLER_211_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07714_ _15409_/Q _07714_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13942__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _08528_/A _08528_/B _08693_/Y vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07940__A _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _07645_/A vssd1 vssd1 vccd1 vccd1 _15443_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07576_ _07576_/A vssd1 vssd1 vccd1 vccd1 _15477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_639 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09315_ _15405_/Q _15389_/Q _09314_/X vssd1 vssd1 vccd1 vccd1 _09320_/B sky130_fd_sc_hd__a21oi_2
XFILLER_139_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14773__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09867__A _15186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _09245_/B _09245_/C _09245_/A vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__o21ai_1
XFILLER_178_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13389__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _09170_/Y _09175_/B _09172_/B vssd1 vssd1 vccd1 vccd1 _09178_/B sky130_fd_sc_hd__o21ai_1
XFILLER_147_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _15008_/Q vssd1 vssd1 vccd1 vccd1 _11687_/A sky130_fd_sc_hd__buf_6
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08059_ _08082_/A _08082_/B _08058_/Y vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__a21oi_1
XFILLER_135_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11070_ _14932_/Q _14998_/Q vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__xor2_2
XFILLER_192_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10021_ _15204_/Q _15105_/Q vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__or2_1
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 x_i_6[12] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 x_i_6[8] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput124 x_i_7[3] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_2
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14013__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput135 x_r_0[13] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input148_A x_r_1[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 x_r_0[9] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput157 x_r_1[4] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__clkbuf_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 x_r_2[14] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__08011__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 x_r_3[0] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__clkbuf_2
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14760_/Y sky130_fd_sc_hd__inv_2
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08489__A1 _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11972_ _11887_/A _11887_/B _11971_/X vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__a21oi_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _13693_/A _13693_/B _13704_/B _13694_/A vssd1 vssd1 vccd1 vccd1 _13718_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _10923_/A _10931_/A vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14691_/Y sky130_fd_sc_hd__inv_2
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13642_ _14971_/Q _13810_/B vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__and2_1
XFILLER_147_1058 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10854_ _10854_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _14919_/D sky130_fd_sc_hd__xor2_2
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11091__B _14935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _15768_/Q _13572_/Y _13571_/A vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__a21o_1
XFILLER_73_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14683__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ _15788_/Q _15722_/Q vssd1 vssd1 vccd1 vccd1 _10786_/B sky130_fd_sc_hd__and2b_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15573_/CLK _15312_/D _14365_/Y vssd1 vssd1 vccd1 vccd1 _15312_/Q sky130_fd_sc_hd__dfrtp_1
X_12524_ _12524_/A _12622_/A vssd1 vssd1 vccd1 vccd1 _15659_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08681__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15243_ _15347_/CLK _15243_/D _14292_/Y vssd1 vssd1 vccd1 vccd1 _15243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12455_ _12455_/A _12455_/B _12455_/C _12455_/D vssd1 vssd1 vccd1 vccd1 _12456_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__10716__A _15283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _15734_/D sky130_fd_sc_hd__xnor2_2
XFILLER_193_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15174_ _15175_/CLK _15174_/D _14218_/Y vssd1 vssd1 vccd1 vccd1 _15174_/Q sky130_fd_sc_hd__dfrtp_1
X_12386_ _12387_/B _12586_/A vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__and2b_1
XFILLER_197_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output367_A output367/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14125_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14125_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _11335_/X _11339_/C vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__and2b_1
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14056_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14056_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13746__B _13746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ _11267_/B _11267_/C _11267_/A vssd1 vssd1 vccd1 vccd1 _11269_/B sky130_fd_sc_hd__a21oi_1
XFILLER_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11547__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ _13091_/A _13007_/B vssd1 vssd1 vccd1 vccd1 _13008_/C sky130_fd_sc_hd__xor2_1
X_10219_ _11400_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _15763_/D sky130_fd_sc_hd__xor2_1
XFILLER_95_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11199_ _15751_/Q _15029_/Q vssd1 vssd1 vccd1 vccd1 _11200_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14858__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater684_A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14958_ _15809_/CLK _14958_/D _13990_/Y vssd1 vssd1 vccd1 vccd1 _14958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _15346_/Q _15330_/Q vssd1 vssd1 vccd1 vccd1 _13909_/X sky130_fd_sc_hd__and2_1
XANTENNA_repeater851_A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14889_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14889_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater949_A input149/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A _15784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07430_ _15548_/Q _07430_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14593__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09100_ _09239_/A _09100_/B vssd1 vssd1 vccd1 vccd1 _15225_/D sky130_fd_sc_hd__xor2_1
XANTENNA__09687__A _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09031_ _09031_/A _09031_/B _13614_/B vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__and3_1
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13937__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09933_ _09932_/A _09932_/B _09990_/B vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__a21o_1
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11457__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _09863_/A _09863_/B _09766_/B vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__a21oi_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _15328_/Q _15344_/Q vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__or2b_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09795_ _09795_/A _09795_/B _09795_/C vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__nor3_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14768__A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08746_ _08631_/X _08633_/A _08745_/X vssd1 vssd1 vccd1 vccd1 _08746_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14918__D _14918_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _12803_/A _12780_/A vssd1 vssd1 vccd1 vccd1 _08677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__A _15750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _15451_/Q input15/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07629_/A sky130_fd_sc_hd__mux2_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ _15485_/Q input49/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07560_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12975__B1 _12976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10570_ _15297_/Q _15264_/Q vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__or2b_1
XFILLER_10_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15749__D _15749_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09227_/A _09227_/B _09228_/X vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__a21o_1
XFILLER_21_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14008__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _12240_/A _12240_/B _12240_/C vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__nand3_1
XFILLER_5_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _12172_/B _12171_/B vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__and2b_1
XFILLER_107_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11122_ _14963_/Q _14897_/Q _11121_/B vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__a21o_1
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13566__B _13567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11053_ _14929_/Q _14995_/Q vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__nand2_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10004_ _15199_/Q _15232_/Q vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__and2_1
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07382__A1 input121/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14678__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14812_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15792_ _15792_/CLK _15792_/D _14872_/Y vssd1 vssd1 vccd1 vccd1 _15792_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__B_N _15751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14743_/Y sky130_fd_sc_hd__inv_2
X_11955_ _11955_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__nand2_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _14962_/Q _14896_/Q vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14674_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14674_/Y sky130_fd_sc_hd__inv_2
X_11886_ _11971_/B _11886_/B vssd1 vssd1 vccd1 vccd1 _11887_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13625_ _13625_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _15099_/D sky130_fd_sc_hd__xor2_1
X_10837_ _10837_/A vssd1 vssd1 vccd1 vccd1 _14913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_780 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13556_ _15765_/Q _13558_/B vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ _10768_/A _10768_/B vssd1 vssd1 vccd1 vccd1 _10769_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output484_A output484/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ _12498_/A _12498_/B _12496_/B _12614_/A _12504_/Y vssd1 vssd1 vccd1 vccd1
+ _12516_/B sky130_fd_sc_hd__a311o_1
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _13416_/A _13180_/C _13259_/A vssd1 vssd1 vccd1 vccd1 _13505_/B sky130_fd_sc_hd__o21ba_1
X_10699_ _10698_/A _10698_/B _11010_/A vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__a21o_1
XFILLER_201_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15226_ _15500_/CLK _15226_/D _14274_/Y vssd1 vssd1 vccd1 vccd1 _15226_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_195_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ _12440_/C _12438_/B _14946_/Q vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__nor3b_1
Xoutput406 output406/A vssd1 vssd1 vccd1 vccd1 y_r_0[3] sky130_fd_sc_hd__buf_2
XFILLER_154_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput417 output417/A vssd1 vssd1 vccd1 vccd1 y_r_1[13] sky130_fd_sc_hd__buf_2
XFILLER_172_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15157_ _15279_/CLK _15157_/D _14201_/Y vssd1 vssd1 vccd1 vccd1 _15157_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput428 _15585_/Q vssd1 vssd1 vccd1 vccd1 y_r_1[8] sky130_fd_sc_hd__buf_2
X_12369_ _12369_/A _12369_/B _12369_/C vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__and3_1
Xoutput439 output439/A vssd1 vssd1 vccd1 vccd1 y_r_2[2] sky130_fd_sc_hd__buf_2
X_14108_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15088_ _15352_/CLK _15088_/D _14128_/Y vssd1 vssd1 vccd1 vccd1 _15088_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__buf_12
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1007 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14588__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__xor2_1
X_09580_ _09580_/A _09795_/A vssd1 vssd1 vccd1 vccd1 _09581_/A sky130_fd_sc_hd__or2_1
XFILLER_167_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ _13319_/A _08531_/B vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__xnor2_2
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08466_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07413_ _07413_/A vssd1 vssd1 vccd1 vccd1 _15561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08393_ _12810_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08396_/C sky130_fd_sc_hd__xor2_1
XFILLER_91_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09014_ _15373_/Q _15357_/Q vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13667__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09916_ _09914_/Y _09916_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11228__B_N _15755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09847_ _15095_/Q _15062_/Q vssd1 vssd1 vccd1 vccd1 _09848_/C sky130_fd_sc_hd__or2b_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14498__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _15155_/D sky130_fd_sc_hd__xnor2_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07604__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08729_ _08728_/A _08728_/B _12627_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08729_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11740_/A _11832_/A _11906_/A vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__and3_1
XFILLER_15_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ _11770_/B _11671_/B vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__xor2_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _13288_/X _13570_/A _13574_/A _13408_/X _13409_/X vssd1 vssd1 vccd1 vccd1
+ _13452_/A sky130_fd_sc_hd__o311ai_4
X_10622_ _10622_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _15001_/D sky130_fd_sc_hd__xor2_1
XFILLER_169_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14390_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14390_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13341_ _13396_/A _13341_/B vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__nand2_2
X_10553_ _10551_/X _10558_/B vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__and2b_1
XFILLER_195_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_956 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13272_ _13272_/A _13272_/B vssd1 vssd1 vccd1 vccd1 _13273_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input76_A x_i_4[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _14903_/D sky130_fd_sc_hd__xor2_1
XFILLER_120_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15011_ _15437_/CLK _15011_/D _14047_/Y vssd1 vssd1 vccd1 vccd1 _15011_/Q sky130_fd_sc_hd__dfrtp_1
X_12223_ _12223_/A _12223_/B _12553_/A _15734_/Q vssd1 vssd1 vccd1 vccd1 _12223_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_154_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13912__A2 _15331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_894 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12154_ _15736_/Q _12154_/B vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11105_ _11105_/A _11105_/B vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__xnor2_1
X_12085_ _12086_/A _12086_/B _12086_/C vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__a21oi_1
XFILLER_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater909 input210/X vssd1 vssd1 vccd1 vccd1 _07850_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11036_ _11311_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14201__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _15775_/CLK _15775_/D _14854_/Y vssd1 vssd1 vccd1 vccd1 _15775_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987_ _13688_/A _13688_/B _12976_/C _12912_/B _12986_/X vssd1 vssd1 vccd1 vccd1
+ _12987_/X sky130_fd_sc_hd__o311a_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14726_/Y sky130_fd_sc_hd__inv_2
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11938_ _12415_/B _11938_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14657_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14657_/Y sky130_fd_sc_hd__inv_2
X_11869_ _12415_/B _11938_/B vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__xor2_2
XFILLER_159_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ _15372_/Q _15356_/Q _13607_/B vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__o21a_1
XFILLER_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14588_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14588_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _15761_/Q _13539_/B vssd1 vssd1 vccd1 vccd1 _13539_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14871__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15209_ _15367_/CLK _15209_/D _14256_/Y vssd1 vssd1 vccd1 vccd1 _15209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput269 output269/A vssd1 vssd1 vccd1 vccd1 y_i_0[2] sky130_fd_sc_hd__buf_2
XFILLER_47_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10623__B _15298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07962_ _10633_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _15004_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _09699_/Y _09701_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1090 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ _07893_/A vssd1 vssd1 vccd1 vccd1 _15321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _09631_/A _09631_/C _09631_/B vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14111__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07424__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09563_ _15435_/Q _15419_/Q vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__nand2_1
XFILLER_71_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09099__A1 _15499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13950__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _14911_/Q vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__buf_6
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _09535_/A _09492_/B _09493_/X vssd1 vssd1 vccd1 vccd1 _15283_/D sky130_fd_sc_hd__a21o_1
XFILLER_211_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08445_ _08464_/A vssd1 vssd1 vccd1 vccd1 _08466_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _13357_/B _08376_/B vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15299__D _15299_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14781__A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_57_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_100_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11629__B _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07585__A1 _07585_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_115_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15762__D _15762_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12910_ _12910_/A _12985_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12912_/A sky130_fd_sc_hd__nand3_2
XFILLER_98_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input130_A x_i_7[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14021__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13890_ _13890_/A _13890_/B vssd1 vssd1 vccd1 vccd1 _15060_/D sky130_fd_sc_hd__xnor2_1
XFILLER_100_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input228_A x_r_6[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12841_ _12841_/A _13669_/B vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__xor2_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15569_/CLK _15560_/D _14627_/Y vssd1 vssd1 vccd1 vccd1 _15560_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12772_ _12772_/A _12772_/B vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__xnor2_4
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14511_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14511_/Y sky130_fd_sc_hd__inv_2
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _12537_/A vssd1 vssd1 vccd1 vccd1 _15581_/D sky130_fd_sc_hd__xnor2_1
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15528_/CLK _15491_/D _14554_/Y vssd1 vssd1 vccd1 vccd1 _15491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A _15754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14442_/Y sky130_fd_sc_hd__inv_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A _12533_/A vssd1 vssd1 vccd1 vccd1 _15580_/D sky130_fd_sc_hd__xor2_1
XFILLER_14_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_759 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10605_ _10532_/Y _10604_/B _10534_/B vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__o21ai_1
X_14373_ _14376_/A vssd1 vssd1 vccd1 vccd1 _14373_/Y sky130_fd_sc_hd__inv_2
X_11585_ _11529_/B _11585_/B vssd1 vssd1 vccd1 vccd1 _11585_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14691__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13324_ _13324_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13325_/B sky130_fd_sc_hd__nor2_1
X_10536_ _10536_/A _10604_/A _10536_/C vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__and3_1
XFILLER_196_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ _13255_/A _13255_/B vssd1 vssd1 vccd1 vccd1 _13257_/B sky130_fd_sc_hd__xor2_1
X_10467_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12206_ _12207_/A _12207_/B _12207_/C vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__a21oi_1
XFILLER_124_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13186_ _13265_/B _13186_/B vssd1 vssd1 vccd1 vccd1 _13187_/B sky130_fd_sc_hd__xnor2_1
X_10398_ _10398_/A vssd1 vssd1 vccd1 vccd1 _14943_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output447_A output447/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ _12186_/A _12137_/B vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09009__B _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater706 _07591_/S vssd1 vssd1 vccd1 vccd1 _07579_/S sky130_fd_sc_hd__buf_4
X_12068_ _12071_/A _12144_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _12074_/A sky130_fd_sc_hd__and3_1
Xrepeater717 _15702_/Q vssd1 vssd1 vccd1 vccd1 output380/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater728 _15680_/Q vssd1 vssd1 vccd1 vccd1 output356/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater597_A _11119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater739 _15660_/Q vssd1 vssd1 vccd1 vccd1 _15813_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08848__B _15446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _11303_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11021_/B sky130_fd_sc_hd__nand2_2
XFILLER_37_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater764_A _15637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14866__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _15758_/CLK _15758_/D _14836_/Y vssd1 vssd1 vccd1 vccd1 _15758_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10635__A1 _15268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater931_A input172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14709_ _14709_/A vssd1 vssd1 vccd1 vccd1 _14709_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15689_ _15689_/CLK _15689_/D _14764_/Y vssd1 vssd1 vccd1 vccd1 _15689_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07500__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11290__A _15786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08230_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__or2_1
XFILLER_20_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ _11480_/A _08201_/B _11617_/A vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08092_ _08109_/A _08108_/A vssd1 vssd1 vccd1 vccd1 _08101_/B sky130_fd_sc_hd__or2_1
XFILLER_134_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14106__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08104__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A1 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13945__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _15369_/Q _15353_/Q vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07945_ _07945_/A vssd1 vssd1 vccd1 vccd1 _15775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07876_ _15329_/Q _07876_/A1 _07892_/S vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__mux2_1
X_09615_ _09615_/A _09615_/B _09809_/A vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__nor3_1
XANTENNA__11184__B _15027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14776__A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09546_ _09545_/A _09545_/B _09775_/A vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__o21a_1
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08774__A _15337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__A2 _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09477_ _15522_/Q _15538_/Q vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__and2b_1
XFILLER_184_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08493__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_737 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08428_ _08429_/A _08429_/B _08427_/Y vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__o21ba_1
XFILLER_34_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _15038_/Q vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__buf_6
XFILLER_20_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11370_ _15751_/Q _15029_/Q _11369_/B vssd1 vssd1 vccd1 vccd1 _11372_/C sky130_fd_sc_hd__a21o_1
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10321_ _10453_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _15781_/D sky130_fd_sc_hd__xnor2_4
XFILLER_137_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14016__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input178_A x_r_2[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _13040_/A _13040_/B vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__or2_1
X_10252_ _10252_/A _10260_/A vssd1 vssd1 vccd1 vccd1 _11411_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10183_ _10183_/A _10854_/A vssd1 vssd1 vccd1 vccd1 _15807_/D sky130_fd_sc_hd__xor2_1
XFILLER_120_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A x_i_2[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _15027_/CLK _14991_/D _14025_/Y vssd1 vssd1 vccd1 vccd1 _14991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13942_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11511__C1 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _15676_/D sky130_fd_sc_hd__xor2_1
XANTENNA__14686__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07730__A1 _07730_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15612_ _15689_/CLK _15612_/D _14683_/Y vssd1 vssd1 vccd1 vccd1 _15612_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ _12921_/A _12822_/Y _12824_/S vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__mux2_1
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08684__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _15561_/CLK _15543_/D _14609_/Y vssd1 vssd1 vccd1 vccd1 _15543_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12755_ _12755_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11706_ _11706_/A _11730_/A vssd1 vssd1 vccd1 vccd1 _11707_/B sky130_fd_sc_hd__xnor2_1
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _15761_/CLK _15474_/D _14536_/Y vssd1 vssd1 vccd1 vccd1 _15474_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _08692_/A _12684_/X _12685_/X vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output397_A output397/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14425_/Y sky130_fd_sc_hd__inv_2
X_11637_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11638_/B sky130_fd_sc_hd__xor2_1
XFILLER_204_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14356_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11568_ _11569_/A _11569_/B _11569_/C vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__a21oi_1
XFILLER_156_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15667__D _15667_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__A1 input236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _13307_/A _13351_/A vssd1 vssd1 vccd1 vccd1 _13308_/C sky130_fd_sc_hd__xnor2_1
XFILLER_115_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10519_ _15257_/Q _15290_/Q vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__nor2_1
X_14287_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14287_/Y sky130_fd_sc_hd__inv_2
X_11499_ _11499_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _11499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13238_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07549__A1 _07549_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _13170_/A _13170_/B _13168_/Y vssd1 vssd1 vccd1 vccd1 _13247_/A sky130_fd_sc_hd__o21bai_2
XFILLER_44_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08859__A _15463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__B _13781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater881_A input245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07730_ _15401_/Q _07730_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater536 _12981_/X vssd1 vssd1 vccd1 vccd1 _15631_/D sky130_fd_sc_hd__clkbuf_2
Xrepeater547 _12525_/X vssd1 vssd1 vccd1 vccd1 _15611_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater558 _11137_/X vssd1 vssd1 vccd1 vccd1 output367/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater569 repeater570/X vssd1 vssd1 vccd1 vccd1 output365/A sky130_fd_sc_hd__buf_4
XFILLER_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07661_ _15435_/Q input255/X _07687_/S vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14596__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _09400_/A _09400_/B vssd1 vssd1 vccd1 vccd1 _15149_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07592_ _07592_/A vssd1 vssd1 vccd1 vccd1 _15469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07702__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ _15409_/Q _15393_/Q vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__xor2_4
XFILLER_209_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _09261_/Y _15489_/Q _09260_/B vssd1 vssd1 vccd1 vccd1 _09265_/B sky130_fd_sc_hd__a21o_1
XFILLER_209_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_193_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _15552_/Q _15572_/Q vssd1 vssd1 vccd1 vccd1 _09195_/A sky130_fd_sc_hd__or2b_1
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08187_/B sky130_fd_sc_hd__xnor2_1
XFILLER_193_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07938__A _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _11458_/A _08290_/B _08074_/C vssd1 vssd1 vccd1 vccd1 _08076_/C sky130_fd_sc_hd__a21oi_1
XFILLER_175_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__A _15336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08977_ _08930_/A _08976_/B _08930_/B vssd1 vssd1 vccd1 vccd1 _15201_/D sky130_fd_sc_hd__a21boi_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07928_ _07928_/A vssd1 vssd1 vccd1 vccd1 _15709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07859_ _07859_/A vssd1 vssd1 vccd1 vccd1 _15338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07712__A1 _07712_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _14957_/Q _14891_/Q vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__or2_1
XFILLER_16_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12738__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _09529_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _15264_/D sky130_fd_sc_hd__xor2_1
XFILLER_43_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _15615_/D sky130_fd_sc_hd__xnor2_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08009__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12471_/A _12471_/B vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__and2_1
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14210_/Y sky130_fd_sc_hd__inv_2
X_11422_ _15082_/Q _15247_/Q vssd1 vssd1 vccd1 vccd1 _11422_/X sky130_fd_sc_hd__and2_1
XFILLER_177_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15190_ _15221_/CLK _15190_/D _14235_/Y vssd1 vssd1 vccd1 vccd1 _15190_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07779__A1 _07779_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14141_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _11353_/A _11353_/B vssd1 vssd1 vccd1 vccd1 _11353_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10304_ _10304_/A _10304_/B vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__nand2_2
XFILLER_3_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14072_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14072_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11284_ _11283_/B _11283_/C _11283_/A vssd1 vssd1 vccd1 vccd1 _11287_/C sky130_fd_sc_hd__a21o_1
XFILLER_193_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13023_ _13023_/A _13023_/B _13023_/C vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__nand3_1
X_10235_ _15077_/Q _15242_/Q vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10166_ _15313_/Q _15148_/Q vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14974_ _15761_/CLK _14974_/D _14007_/Y vssd1 vssd1 vccd1 vccd1 _14974_/Q sky130_fd_sc_hd__dfrtp_2
X_10097_ _15217_/Q _15118_/Q vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__xnor2_2
X_13925_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13925_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12929__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_795 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13856_ _13859_/B _13856_/B vssd1 vssd1 vccd1 vccd1 _15672_/D sky130_fd_sc_hd__nor2_1
XFILLER_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07522__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _12807_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _12807_/Y sky130_fd_sc_hd__nor2_1
X_13787_ _14984_/Q _13867_/B vssd1 vssd1 vccd1 vccd1 _13788_/B sky130_fd_sc_hd__or2_1
XFILLER_204_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10999_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__and3_1
XFILLER_128_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12738_ _13145_/A _12970_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__and3_1
X_15526_ _15528_/CLK _15526_/D _14591_/Y vssd1 vssd1 vccd1 vccd1 _15526_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15457_ _15700_/CLK _15457_/D _14518_/Y vssd1 vssd1 vccd1 vccd1 _15457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12669_ _12803_/A _08499_/C _12668_/Y vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater727_A _15685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14408_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14408_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _15411_/CLK _15388_/D _14446_/Y vssd1 vssd1 vccd1 vccd1 _15388_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14339_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08900_ _08900_/A _08900_/B _08959_/B vssd1 vssd1 vccd1 vccd1 _08900_/X sky130_fd_sc_hd__and3_1
XFILLER_83_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__nand2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08836_/A vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__or2_1
XFILLER_111_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08762_ _15333_/Q _08763_/B _13874_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__a21oi_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07713_ _07713_/A vssd1 vssd1 vccd1 vccd1 _15410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08693_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08693_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07644_ _15443_/Q _07644_/A1 _07644_/S vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07940__B _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07432__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07575_ _15477_/Q _07575_/A1 _07575_/S vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09314_ _15405_/Q _15389_/Q _09310_/B vssd1 vssd1 vccd1 vccd1 _09314_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09245_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__or3_1
XFILLER_181_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12574__A _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ _15569_/Q _15549_/Q vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__xnor2_1
XFILLER_147_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08127_ _15010_/Q vssd1 vssd1 vccd1 vccd1 _11832_/A sky130_fd_sc_hd__buf_6
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07630__A0 _15450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _08058_/A _08058_/B vssd1 vssd1 vccd1 vccd1 _08058_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_747 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08499__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ _10020_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _14972_/D sky130_fd_sc_hd__xnor2_2
Xinput103 x_i_6[13] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput114 x_i_6[9] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 x_i_7[4] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__buf_4
XFILLER_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 x_r_0[14] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput147 x_r_1[0] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput158 x_r_1[5] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08011__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 x_r_2[15] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11971_ _11886_/B _11971_/B vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__and2b_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08489__A2 _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_710 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13710_ _13703_/A _13700_/X _13703_/B vssd1 vssd1 vccd1 vccd1 _13718_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input210_A x_r_4[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _14898_/Q _14964_/Q vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__or2b_1
X_14690_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14690_/Y sky130_fd_sc_hd__inv_2
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13641_ _13641_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _15693_/D sky130_fd_sc_hd__xnor2_1
X_10853_ _10852_/A _10852_/B _10175_/B vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13572_/A vssd1 vssd1 vccd1 vccd1 _13572_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10784_ _15722_/Q _15788_/Q vssd1 vssd1 vccd1 vccd1 _10786_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08962__A _15471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15573_/CLK _15311_/D _14364_/Y vssd1 vssd1 vccd1 vccd1 _15311_/Q sky130_fd_sc_hd__dfrtp_2
X_12523_ _12523_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12622_/A sky130_fd_sc_hd__xnor2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_858 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15347_/CLK _15242_/D _14291_/Y vssd1 vssd1 vccd1 vccd1 _15242_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12454_ _12454_/A _12454_/B _12455_/C vssd1 vssd1 vccd1 vccd1 _12456_/C sky130_fd_sc_hd__or3b_1
XANTENNA__13299__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _10230_/A _11404_/B _10230_/B vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__a21boi_2
XFILLER_172_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15173_ _15175_/CLK _15173_/D _14217_/Y vssd1 vssd1 vccd1 vccd1 _15173_/Q sky130_fd_sc_hd__dfrtp_1
X_12385_ _12383_/Y _12385_/B vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__and2b_1
XFILLER_193_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14124_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ _11335_/B _11335_/C _11335_/A vssd1 vssd1 vccd1 vccd1 _11339_/C sky130_fd_sc_hd__a21o_1
XFILLER_180_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output262_A output262/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14055_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14055_/Y sky130_fd_sc_hd__inv_2
X_11267_ _11267_/A _11267_/B _11267_/C vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__and3_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14204__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13006_ _13006_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__nand2_1
X_10218_ _15073_/Q _10217_/Y _10213_/B vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08202__A _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11198_ _15751_/Q _15029_/Q vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__or2_1
XANTENNA_output527_A output527/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10150_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14957_ _15809_/CLK _14957_/D _13989_/Y vssd1 vssd1 vccd1 vccd1 _14957_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater677_A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13908_/A _13908_/B vssd1 vssd1 vccd1 vccd1 _15066_/D sky130_fd_sc_hd__xor2_1
XFILLER_169_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14888_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14888_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12378__B _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater844_A repeater845/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13839_ _13838_/A _13838_/C _13838_/B vssd1 vssd1 vccd1 vccd1 _13842_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14874__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__A _15467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15509_ _15509_/CLK _15509_/D _14573_/Y vssd1 vssd1 vccd1 vccd1 _15509_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_206_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ _09030_/A _09038_/A vssd1 vssd1 vccd1 vccd1 _13614_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07860__A0 _15337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__B _15299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09932_ _09932_/A _09932_/B _09990_/B vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__and3_1
XFILLER_131_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14114__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _15757_/D sky130_fd_sc_hd__xor2_1
XFILLER_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13953__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08814_/A vssd1 vssd1 vccd1 vccd1 _15079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09580_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09795_/C sky130_fd_sc_hd__and2b_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08715_/Y _08717_/X _08713_/Y vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__a21bo_1
XFILLER_45_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11473__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__A0 _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _12970_/A _12803_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__and3_1
XFILLER_27_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__B _15028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ _07627_/A vssd1 vssd1 vccd1 vccd1 _15452_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14784__A _14784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07558_ _07558_/A vssd1 vssd1 vccd1 vccd1 _15486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14934__D _14934_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07489_ _07489_/A vssd1 vssd1 vccd1 vccd1 _15520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _15496_/Q _15480_/Q vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__and2b_1
XFILLER_42_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12727__A1 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _09153_/Y _09157_/B _09155_/B vssd1 vssd1 vccd1 vccd1 _09160_/B sky130_fd_sc_hd__o21ai_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12170_ _12238_/A _12109_/Y _12111_/A _12169_/Y vssd1 vssd1 vccd1 vccd1 _12171_/B
+ sky130_fd_sc_hd__o31ai_1
X_11121_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_190_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input160_A x_r_1[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input258_A x_r_7[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14024__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09118__A _15488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _14929_/Q _14995_/Q vssd1 vssd1 vccd1 vccd1 _11052_/Y sky130_fd_sc_hd__nor2_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _14935_/D sky130_fd_sc_hd__xor2_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input21_A x_i_1[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14811_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14811_/Y sky130_fd_sc_hd__inv_2
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _15791_/CLK _15791_/D _14871_/Y vssd1 vssd1 vccd1 vccd1 _15791_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_946 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11383__A _15755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ _11954_/A vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__inv_2
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14753_/A sky130_fd_sc_hd__buf_6
XFILLER_45_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _10905_/A vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14673_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14673_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11885_ _11960_/A _11668_/C _12055_/A vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14694__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13624_ _13622_/A _13622_/B _13623_/X vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__a21o_1
X_10836_ _10836_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10837_/A sky130_fd_sc_hd__and2_1
XFILLER_16_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13555_ _13555_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _15601_/D sky130_fd_sc_hd__xnor2_1
XFILLER_201_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10767_ _15718_/Q _15784_/Q _10763_/B vssd1 vssd1 vccd1 vccd1 _10768_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _12614_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13103__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13486_ _13473_/A _13473_/B _13471_/A vssd1 vssd1 vccd1 vccd1 _13505_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ _10698_/A _10698_/B _11010_/A vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__and3_1
XFILLER_139_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output477_A _11269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15225_ _15500_/CLK _15225_/D _14273_/Y vssd1 vssd1 vccd1 vccd1 _15225_/Q sky130_fd_sc_hd__dfrtp_1
X_12437_ _12437_/A vssd1 vssd1 vccd1 vccd1 _15651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput407 output407/A vssd1 vssd1 vccd1 vccd1 y_r_0[4] sky130_fd_sc_hd__buf_2
X_15156_ _15279_/CLK _15156_/D _14200_/Y vssd1 vssd1 vccd1 vccd1 _15156_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput418 _15591_/Q vssd1 vssd1 vccd1 vccd1 y_r_1[14] sky130_fd_sc_hd__buf_2
X_12368_ _14941_/Q vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__inv_2
Xoutput429 output429/A vssd1 vssd1 vccd1 vccd1 y_r_1[9] sky130_fd_sc_hd__buf_2
XFILLER_181_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14107_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11319_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__and3_1
XFILLER_141_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _15352_/CLK _15087_/D _14127_/Y vssd1 vssd1 vccd1 vccd1 _15087_/Q sky130_fd_sc_hd__dfrtp_1
X_12299_ _15738_/Q vssd1 vssd1 vccd1 vccd1 _12299_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14038_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__buf_12
XFILLER_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14869__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater794_A _15595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater961_A input133/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ _08530_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ _08592_/A _08594_/A vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__and2b_1
XFILLER_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07412_ _15561_/Q _07412_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07413_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08392_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08392_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07710__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__B _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10637__A _15269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14109__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _15373_/Q _15357_/Q vssd1 vssd1 vccd1 vccd1 _09013_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12709__A1 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13948__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13382__A1 _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A _15251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09915_ _15193_/Q _15226_/Q vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14779__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _15431_/Q _15415_/Q _09776_/X vssd1 vssd1 vccd1 vccd1 _09778_/B sky130_fd_sc_hd__a21o_1
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _08728_/A _08728_/B _12627_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08728_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08659_ _08427_/A _08427_/B _08658_/Y vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__a21oi_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11764_/A _11445_/B _11876_/A vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__mux2_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ _10619_/A _10619_/B _10620_/X vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14019__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13340_ _13340_/A _13340_/B _13340_/C vssd1 vssd1 vccd1 vccd1 _13341_/B sky130_fd_sc_hd__nand3_1
XFILLER_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10552_ _10551_/A _10551_/B _10609_/B vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__a21o_1
XFILLER_183_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08017__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13270_/A _13270_/B _13270_/C vssd1 vssd1 vccd1 vccd1 _13272_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ _10482_/A _10482_/B _10367_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15010_ _15437_/CLK _15010_/D _14046_/Y vssd1 vssd1 vccd1 vccd1 _15010_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12222_ _12560_/A _12220_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__or2b_1
XFILLER_120_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input69_A x_i_4[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12153_ _15736_/Q _12154_/B vssd1 vssd1 vccd1 vccd1 _12220_/A sky130_fd_sc_hd__and2_1
XFILLER_190_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _11104_/A _11352_/A vssd1 vssd1 vccd1 vccd1 _11104_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_155_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11097__B _15002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ _12141_/B _12084_/B vssd1 vssd1 vccd1 vccd1 _12086_/C sky130_fd_sc_hd__or2_1
XFILLER_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14689__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11035_ _11029_/A _11031_/B _11029_/B vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__a21boi_1
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12884__B1 _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _13677_/A _12986_/B vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__or2_1
X_15774_ _15774_/CLK _15774_/D _14853_/Y vssd1 vssd1 vccd1 vccd1 _15774_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14725_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14725_/Y sky130_fd_sc_hd__inv_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _12426_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__xnor2_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ _11868_/A _11868_/B vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__xor2_2
X_14656_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14656_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07530__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10819_ _10817_/A _10817_/B _10818_/X vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__a21o_1
X_13607_ _13607_/A _13607_/B vssd1 vssd1 vccd1 vccd1 _15093_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_repeater542_A _10958_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11799_ _11799_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11811_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14587_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14587_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13538_ _15761_/Q _13539_/B vssd1 vssd1 vccd1 vccd1 _13538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09280__A2 _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13469_ _13470_/A _13470_/B _13470_/C vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater807_A _15582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12672__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ _15367_/CLK _15208_/D _14255_/Y vssd1 vssd1 vccd1 vccd1 _15208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15139_ _15406_/CLK _15139_/D _14182_/Y vssd1 vssd1 vccd1 vccd1 _15139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput259 output259/A vssd1 vssd1 vccd1 vccd1 finish sky130_fd_sc_hd__buf_2
XFILLER_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ _15152_/Q _15251_/Q vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14599__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _15057_/Q _15090_/Q vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07892_ _15321_/Q _07892_/A1 _07892_/S vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09633_/A sky130_fd_sc_hd__and3_1
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11735__B _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09562_ _15435_/Q _15419_/Q vssd1 vssd1 vccd1 vccd1 _09562_/Y sky130_fd_sc_hd__nor2_1
X_08513_ _12970_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09493_ _15540_/Q _15524_/Q vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ _08444_/A _08466_/C vssd1 vssd1 vccd1 vccd1 _08587_/A sky130_fd_sc_hd__xnor2_1
XFILLER_63_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08375_ _08371_/A _08371_/B _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08408_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_11_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07806__A0 _15364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11198__A _15751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13107__A1 _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14302__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09829_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _15747_/D sky130_fd_sc_hd__xor2_2
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12840_ _13677_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13669_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_input123_A x_i_7[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08298__B1 _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _12772_/B sky130_fd_sc_hd__nand2_2
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _15730_/Q _11725_/B vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__xnor2_4
X_14510_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14510_/Y sky130_fd_sc_hd__inv_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15500_/CLK _15490_/D _14553_/Y vssd1 vssd1 vccd1 vccd1 _15490_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11380__B _15032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11653_ _15729_/Q _12534_/B vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__xnor2_2
X_14441_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14460_/A sky130_fd_sc_hd__buf_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10604_ _10604_/A _10604_/B vssd1 vssd1 vccd1 vccd1 _14995_/D sky130_fd_sc_hd__xnor2_1
X_14372_ _14376_/A vssd1 vssd1 vccd1 vccd1 _14372_/Y sky130_fd_sc_hd__inv_2
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13323_ _13438_/A _13390_/A _13381_/B vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__and3b_1
XFILLER_11_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ _15291_/Q _15258_/Q vssd1 vssd1 vccd1 vccd1 _10536_/C sky130_fd_sc_hd__or2b_1
XFILLER_155_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13254_ _13366_/A _12927_/B _13300_/A vssd1 vssd1 vccd1 vccd1 _13255_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10466_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _14897_/D sky130_fd_sc_hd__xor2_1
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12205_ _12256_/B _12205_/B vssd1 vssd1 vccd1 vccd1 _12207_/C sky130_fd_sc_hd__nand2_1
XFILLER_170_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13253_/B _12888_/C _13357_/B vssd1 vssd1 vccd1 vccd1 _13186_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ _10397_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__and2_1
XFILLER_151_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12136_ _12193_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12137_/B sky130_fd_sc_hd__and2_1
XFILLER_111_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output342_A output342/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11836__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ _12204_/A vssd1 vssd1 vccd1 vccd1 _12071_/A sky130_fd_sc_hd__inv_2
XANTENNA__14212__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater707 _07575_/S vssd1 vssd1 vccd1 vccd1 _07591_/S sky130_fd_sc_hd__buf_6
Xrepeater718 _15701_/Q vssd1 vssd1 vccd1 vccd1 output395/A sky130_fd_sc_hd__clkbuf_2
Xrepeater729 _15679_/Q vssd1 vssd1 vccd1 vccd1 output355/A sky130_fd_sc_hd__clkbuf_2
X_11018_ _14922_/Q _14988_/Q vssd1 vssd1 vccd1 vccd1 _11019_/B sky130_fd_sc_hd__or2b_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13770__B _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15758_/CLK _15757_/D _14835_/Y vssd1 vssd1 vccd1 vccd1 _15757_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater757_A _15644_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _13048_/B _12969_/B vssd1 vssd1 vccd1 vccd1 _12970_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12667__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14708_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15688_ _15688_/CLK _15688_/D _14763_/Y vssd1 vssd1 vccd1 vccd1 _15688_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater924_A input185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14639_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14882__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08160_ _11687_/A _11491_/A vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__xor2_1
XFILLER_165_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08091_ _11898_/A _08097_/B vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__nand2_1
XFILLER_162_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08104__B _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08993_ _15369_/Q _15353_/Q vssd1 vssd1 vccd1 vccd1 _08993_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07943__B _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _10295_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__and2_1
XFILLER_69_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10650__A _15272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14122__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07435__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07875_ _07875_/A vssd1 vssd1 vccd1 vccd1 _15330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13961__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ _15443_/Q _15427_/Q vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09545_ _09545_/A _09545_/B _09775_/A vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__nor3_1
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_129_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08774__B _15321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _09476_/A vssd1 vssd1 vccd1 vccd1 _15279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12296__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14792__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08358_ _15040_/Q vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__buf_6
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14942__D _14942_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _08289_/A _08289_/B vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__xor2_2
XFILLER_192_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _10314_/A _10316_/B _10314_/B vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__13201__A _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _15244_/Q _15079_/Q vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__or2b_1
XFILLER_182_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__nor2_2
XFILLER_160_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input240_A x_r_6[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ _15119_/CLK _14990_/D _14024_/Y vssd1 vssd1 vccd1 vccd1 _14990_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14032__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09126__A _15505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13941_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13871__A _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13872_ _13868_/A _13870_/X _13868_/B _13871_/X vssd1 vssd1 vccd1 vccd1 _13873_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_46_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15611_ _15706_/CLK _15611_/D _14681_/Y vssd1 vssd1 vccd1 vccd1 _15611_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12823_ _12945_/A vssd1 vssd1 vccd1 vccd1 _12824_/S sky130_fd_sc_hd__inv_2
XFILLER_15_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08684__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ _15542_/CLK _15542_/D _14608_/Y vssd1 vssd1 vccd1 vccd1 _15542_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12755_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11705_ _11705_/A _11733_/A vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__xor2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07494__A1 _07494_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__and2_1
X_15473_ _15511_/CLK _15473_/D _14535_/Y vssd1 vssd1 vccd1 vccd1 _15473_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _11558_/A _11558_/B _11635_/Y vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__a21o_1
X_14424_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14424_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output292_A output292/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11567_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11569_/C sky130_fd_sc_hd__xnor2_1
XFILLER_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14355_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14355_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14207__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10518_ _10598_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _15025_/D sky130_fd_sc_hd__xor2_1
X_13306_ _13255_/A _13255_/B _13258_/B vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__a21oi_1
XFILLER_171_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14286_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14286_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08205__A _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11498_ _11499_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _11498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13333_/B sky130_fd_sc_hd__and2_1
X_10449_ _15123_/Q _10448_/Y _10447_/B vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _13220_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13168_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15683__D _15683_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12119_/A _12119_/B _12119_/C vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__or3_1
X_13099_ _13100_/A _13100_/B _13100_/C vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09036__A _15376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater537 _11350_/X vssd1 vssd1 vccd1 vccd1 output334/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14877__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater548 _11344_/X vssd1 vssd1 vccd1 vccd1 output331/A sky130_fd_sc_hd__clkbuf_2
Xrepeater559 _10940_/X vssd1 vssd1 vccd1 vccd1 _10941_/A sky130_fd_sc_hd__buf_2
XANTENNA__13781__A _13781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _07660_/A vssd1 vssd1 vccd1 vccd1 _15436_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_56_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15809_ _15809_/CLK _15809_/D _14889_/Y vssd1 vssd1 vccd1 vccd1 _15809_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07591_ _15469_/Q _07591_/A1 _07591_/S vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09330_ _09328_/A _09386_/B _09329_/X vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__a21o_2
XFILLER_206_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _15505_/Q vssd1 vssd1 vccd1 vccd1 _09261_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ _08292_/B _08218_/B _08219_/B _08211_/X vssd1 vssd1 vccd1 vccd1 _08215_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ _15571_/Q _15551_/Q _09191_/B vssd1 vssd1 vccd1 vccd1 _09196_/A sky130_fd_sc_hd__a21o_1
XFILLER_140_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_114_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _11707_/A _11617_/A vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10645__A _15271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14117__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08074_ _11458_/A _15792_/Q _08074_/C vssd1 vssd1 vccd1 vccd1 _08094_/A sky130_fd_sc_hd__and3_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13956__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12860__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11741__A0 _11842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11476__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10380__A _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08976_ _08976_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _15200_/D sky130_fd_sc_hd__xnor2_1
XFILLER_88_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07927_ _09686_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__and2_1
XFILLER_116_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07858_ _15338_/Q input206/X _07900_/S vssd1 vssd1 vccd1 vccd1 _07859_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _15372_/Q _07789_/A1 _07791_/S vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09526_/A _09526_/B _09527_/X vssd1 vssd1 vccd1 vccd1 _09529_/B sky130_fd_sc_hd__a21o_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09459_/A _09459_/B _09518_/B vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__and3_1
XFILLER_196_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08009__B _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ _14949_/Q _12484_/B _12475_/C vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__nand3b_1
XFILLER_71_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11421_ _11421_/A _11421_/B vssd1 vssd1 vccd1 vccd1 _15739_/D sky130_fd_sc_hd__xor2_2
XANTENNA_input190_A x_r_3[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14027__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14140_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14140_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11352_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11352_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_180_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ _15122_/Q _15155_/Q vssd1 vssd1 vccd1 vccd1 _10304_/B sky130_fd_sc_hd__nand2_1
X_14071_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14071_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _11283_/A _11283_/B _11283_/C vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__and3_1
XFILLER_3_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13022_ _13022_/A _13022_/B _13022_/C _13022_/D vssd1 vssd1 vccd1 vccd1 _13023_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA_input51_A x_i_3[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10234_ _11404_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10239_/A sky130_fd_sc_hd__nand2_1
XFILLER_193_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07400__A1 _07400_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__A _15756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _15148_/Q _15313_/Q vssd1 vssd1 vccd1 vccd1 _10167_/A sky130_fd_sc_hd__and2b_1
XFILLER_79_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14973_ _15493_/CLK _14973_/D _14006_/Y vssd1 vssd1 vccd1 vccd1 _14973_/Q sky130_fd_sc_hd__dfrtp_1
X_10096_ _10094_/A _10432_/A _10095_/Y vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__14697__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_590 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13924_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13924_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12929__B _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13855_ _13848_/A _13848_/B _13849_/X _13767_/B vssd1 vssd1 vccd1 vccd1 _13856_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA_output305_A output305/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13106__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ _12804_/Y _13056_/B vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__and2b_1
X_10998_ _15177_/Q _15276_/Q vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__or2b_1
X_13786_ _14984_/Q _13867_/B vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__A1 _07467_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15525_ _15525_/CLK _15525_/D _14590_/Y vssd1 vssd1 vccd1 vccd1 _15525_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12737_ _12871_/A _12803_/A _12780_/A vssd1 vssd1 vccd1 vccd1 _12781_/A sky130_fd_sc_hd__and3b_1
XFILLER_96_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12945__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15456_ _15571_/CLK _15456_/D _14517_/Y vssd1 vssd1 vccd1 vccd1 _15456_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ _12871_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _12668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14407_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14407_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11619_ _11562_/A _11562_/B _11618_/X vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_repeater622_A _10743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15387_ _15392_/CLK _15387_/D _14445_/Y vssd1 vssd1 vccd1 vccd1 _15387_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12599_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _15685_/D sky130_fd_sc_hd__xnor2_1
XFILLER_128_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14338_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14269_ _14269_/A vssd1 vssd1 vccd1 vccd1 _14269_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _15346_/Q _15330_/Q vssd1 vssd1 vccd1 vccd1 _08836_/A sky130_fd_sc_hd__and2b_1
XFILLER_140_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08766_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__or2_1
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07712_ _15410_/Q _07712_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08692_ _08692_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__14400__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07643_ _07643_/A vssd1 vssd1 vccd1 vccd1 _15444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07574_ _07574_/A vssd1 vssd1 vccd1 vccd1 _15478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09313_ _09320_/A _09321_/A vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__or2_1
XFILLER_62_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15732_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09244_ _15501_/Q _15485_/Q vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__and2b_1
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15588__D _15588_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09175_ _09648_/A _09175_/B vssd1 vssd1 vccd1 vccd1 _15291_/D sky130_fd_sc_hd__xor2_1
XFILLER_31_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08126_ _15007_/Q vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__buf_4
XFILLER_147_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08057_ _08290_/B _08057_/B vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07630__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08499__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 x_i_6[14] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__clkbuf_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput115 x_i_7[0] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_2
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput126 x_i_7[5] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput137 x_r_0[15] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__clkbuf_2
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 x_r_1[10] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_4
XFILLER_103_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput159 x_r_1[6] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08959_ _08959_/A _08959_/B _08959_/C vssd1 vssd1 vccd1 vccd1 _08961_/A sky130_fd_sc_hd__nor3_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11970_ _12030_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__xnor2_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14310__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07697__A1 input189/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _14964_/Q _14898_/Q vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__or2b_1
XFILLER_17_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater890 input234/X vssd1 vssd1 vccd1 vccd1 _07801_/A1 sky130_fd_sc_hd__buf_4
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input203_A x_r_4[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _10852_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _14918_/D sky130_fd_sc_hd__xor2_2
X_13640_ _13810_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13809_/B sky130_fd_sc_hd__xnor2_4
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07449__A1 _07449_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10783_ _15721_/Q _15787_/Q vssd1 vssd1 vccd1 vccd1 _10787_/B sky130_fd_sc_hd__nand2_1
X_13571_ _13571_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _15604_/D sky130_fd_sc_hd__nor2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15383_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08962__B _15455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15573_/CLK _15310_/D _14363_/Y vssd1 vssd1 vccd1 vccd1 _15310_/Q sky130_fd_sc_hd__dfrtp_1
X_12522_ _14954_/Q _12522_/B vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__xor2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input99_A x_i_6[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _15347_/CLK _15241_/D _14290_/Y vssd1 vssd1 vccd1 vccd1 _15241_/Q sky130_fd_sc_hd__dfrtp_1
X_12453_ _12416_/A _12455_/A _12430_/C vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13299__C _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08949__A1 _15466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _15733_/D sky130_fd_sc_hd__xnor2_2
X_12384_ _12384_/A _12391_/C _12389_/C vssd1 vssd1 vccd1 vccd1 _12385_/B sky130_fd_sc_hd__nand3_1
X_15172_ _15433_/CLK _15172_/D _14216_/Y vssd1 vssd1 vccd1 vccd1 _15172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14123_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14123_/Y sky130_fd_sc_hd__inv_2
X_11335_ _11335_/A _11335_/B _11335_/C vssd1 vssd1 vccd1 vccd1 _11335_/X sky130_fd_sc_hd__and3_1
XFILLER_193_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14054_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__inv_2
X_11266_ _15780_/Q _15714_/Q vssd1 vssd1 vccd1 vccd1 _11267_/C sky130_fd_sc_hd__or2b_1
XFILLER_122_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13005_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__xnor2_1
X_10217_ _15238_/Q vssd1 vssd1 vccd1 vccd1 _10217_/Y sky130_fd_sc_hd__inv_2
X_11197_ _11197_/A _11197_/B vssd1 vssd1 vccd1 vccd1 _11197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_451 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _15144_/Q _15309_/Q _10144_/B vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output422_A _15579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14956_ _15809_/CLK _14956_/D _13988_/Y vssd1 vssd1 vccd1 vccd1 _14956_/Q sky130_fd_sc_hd__dfrtp_1
X_10079_ _10079_/A _10079_/B _10428_/A vssd1 vssd1 vccd1 vccd1 _10079_/X sky130_fd_sc_hd__and3_1
XANTENNA__14220__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13907_ _13905_/A _13905_/B _13906_/X vssd1 vssd1 vccd1 vccd1 _13908_/B sky130_fd_sc_hd__a21o_1
XFILLER_208_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14887_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _13838_/A _13838_/B _13838_/C vssd1 vssd1 vccd1 vccd1 _13840_/A sky130_fd_sc_hd__nor3_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _13769_/A _13769_/B vssd1 vssd1 vccd1 vccd1 _13783_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12675__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15799_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08872__B _15451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15508_ _15508_/CLK _15508_/D _14572_/Y vssd1 vssd1 vccd1 vccd1 _15508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _15439_/CLK _15439_/D _14499_/Y vssd1 vssd1 vccd1 vccd1 _15439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07860__A1 input205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07612__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07708__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _09931_/A _09939_/A vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09861_/A _09861_/B _09759_/B vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__a21o_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _08811_/X _08818_/B vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__and2b_1
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _15161_/D sky130_fd_sc_hd__xnor2_1
XFILLER_133_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09117__A1 _15503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _08714_/X _08719_/X _08720_/X _08743_/X vssd1 vssd1 vccd1 vccd1 _08744_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14130__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11473__B _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08675_ _12780_/A _08675_/B vssd1 vssd1 vccd1 vccd1 _08680_/A sky130_fd_sc_hd__nor2_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07626_ _15452_/Q input16/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07627_/A sky130_fd_sc_hd__mux2_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ _15486_/Q input50/X _07591_/S vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15588_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07488_ _15520_/Q input21/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10986__A1 _15273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09227_ _09227_/A _09227_/B vssd1 vssd1 vccd1 vccd1 _15237_/D sky130_fd_sc_hd__xor2_2
XFILLER_10_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ _15565_/Q _15545_/Q vssd1 vssd1 vccd1 vccd1 _09639_/A sky130_fd_sc_hd__xnor2_2
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08304_/B sky130_fd_sc_hd__xor2_1
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14950__D _14950_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09089_ _15497_/Q _15481_/Q _09085_/B vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14305__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ _10906_/Y _11119_/B _10908_/B vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__o21ai_4
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A_N _15462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11051_ _11325_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11051_/Y sky130_fd_sc_hd__xnor2_2
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input153_A x_r_1[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10002_ _10000_/A _10000_/B _10001_/X vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__a21o_1
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15781__D _15781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14810_/Y sky130_fd_sc_hd__inv_2
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14040__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _15790_/CLK _15790_/D _14870_/Y vssd1 vssd1 vccd1 vccd1 _15790_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A x_i_0[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__B _15033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _14741_/A vssd1 vssd1 vccd1 vccd1 _14741_/Y sky130_fd_sc_hd__inv_2
X_11953_ _11896_/B _11953_/B vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__and2b_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ _10904_/A _10910_/A vssd1 vssd1 vccd1 vccd1 _10905_/A sky130_fd_sc_hd__and2_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14672_/Y sky130_fd_sc_hd__inv_2
X_11884_ _12122_/A vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__inv_2
XFILLER_45_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_13623_ _15377_/Q _15361_/Q vssd1 vssd1 vccd1 vccd1 _13623_/X sky130_fd_sc_hd__and2_1
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10835_ _10834_/B _10834_/C _10834_/A vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__o21ai_1
XFILLER_186_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13554_ _13551_/A _13552_/A _13551_/B _13066_/B _13553_/Y vssd1 vssd1 vccd1 vccd1
+ _13560_/B sky130_fd_sc_hd__o32a_1
XFILLER_185_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10766_ _10766_/A _11287_/A vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12498_/A _12498_/B _12496_/B _12504_/Y vssd1 vssd1 vccd1 vccd1 _12506_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13103__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07842__A1 _07842_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _10697_/A _10697_/B vssd1 vssd1 vccd1 vccd1 _11010_/A sky130_fd_sc_hd__nor2_1
X_13485_ _13475_/A _13483_/Y _13484_/X vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__a21o_1
XFILLER_12_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _15483_/CLK _15224_/D _14272_/Y vssd1 vssd1 vccd1 vccd1 _15224_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12436_ _12478_/A _12436_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__and2b_1
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output372_A _11109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11839__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15155_ _15279_/CLK _15155_/D _14198_/Y vssd1 vssd1 vccd1 vccd1 _15155_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput408 output408/A vssd1 vssd1 vccd1 vccd1 y_r_0[5] sky130_fd_sc_hd__buf_2
X_12367_ _12364_/A _12578_/A _12366_/Y vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__a21o_1
Xoutput419 output419/A vssd1 vssd1 vccd1 vccd1 y_r_1[15] sky130_fd_sc_hd__buf_2
XANTENNA__14215__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07528__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14106_/Y sky130_fd_sc_hd__inv_2
X_11318_ _14992_/Q _14926_/Q vssd1 vssd1 vccd1 vccd1 _11319_/C sky130_fd_sc_hd__or2b_1
X_12298_ _12298_/A _12567_/A vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__nor2_1
X_15086_ _15367_/CLK _15086_/D _14126_/Y vssd1 vssd1 vccd1 vccd1 _15086_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11249_ _15775_/Q _11248_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _11251_/C sky130_fd_sc_hd__a21o_1
X_14037_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14037_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater787_A repeater788/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14939_ _15727_/CLK _14939_/D _13970_/Y vssd1 vssd1 vccd1 vccd1 _14939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater954_A input142/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14885__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__nor2_1
XFILLER_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07530__A0 _15499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07411_ _07411_/A vssd1 vssd1 vccd1 vccd1 _15562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ _08391_/A _08391_/B vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13603__B1 _13602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15027_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_211_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11740__C _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ _13607_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _15109_/D sky130_fd_sc_hd__xor2_1
XFILLER_176_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12709__A2 _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14125__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09219__A _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13964__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09914_ _15193_/Q _15226_/Q vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A x_i_0[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13683__B _13824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _15751_/D sky130_fd_sc_hd__xor2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09776_ _15431_/Q _15415_/Q _09775_/B vssd1 vssd1 vccd1 vccd1 _09776_/X sky130_fd_sc_hd__o21a_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08727_ _12654_/A _12688_/A _08726_/Y vssd1 vssd1 vccd1 vccd1 _08727_/X sky130_fd_sc_hd__a21o_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11448__A2 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14795__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08658_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08658_/Y sky130_fd_sc_hd__nor2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07609_/A vssd1 vssd1 vccd1 vccd1 _15461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14945__D _14945_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08589_/A _08589_/B vssd1 vssd1 vccd1 vccd1 _08713_/A sky130_fd_sc_hd__xnor2_2
XFILLER_186_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10620_ _15264_/Q _15297_/Q vssd1 vssd1 vccd1 vccd1 _10620_/X sky130_fd_sc_hd__and2_1
XFILLER_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__A1 input175/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ _10551_/A _10551_/B _10609_/B vssd1 vssd1 vccd1 vccd1 _10551_/X sky130_fd_sc_hd__and3_1
XANTENNA__08017__B _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _14902_/D sky130_fd_sc_hd__xor2_1
X_13270_ _13270_/A _13270_/B _13270_/C vssd1 vssd1 vccd1 vccd1 _13272_/A sky130_fd_sc_hd__and3_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15776__D _15776_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12221_ _12560_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_68_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14035__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12152_ _12152_/A _12456_/A vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ _14937_/Q _15003_/Q vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__xnor2_4
XFILLER_123_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08968__A _08968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _11032_/Y _11034_/B vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__and2b_1
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08179__S _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/CLK _15773_/D _14852_/Y vssd1 vssd1 vccd1 vccd1 _15773_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_17_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12985_ _13020_/B _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _13688_/B sky130_fd_sc_hd__and3b_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14724_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14724_/Y sky130_fd_sc_hd__inv_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__xor2_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14655_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14655_/Y sky130_fd_sc_hd__inv_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11868_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _09003_/Y _13605_/B _09005_/B vssd1 vssd1 vccd1 vccd1 _13607_/B sky130_fd_sc_hd__o21ai_1
X_10818_ _15304_/Q _15139_/Q vssd1 vssd1 vccd1 vccd1 _10818_/X sky130_fd_sc_hd__and2b_1
XFILLER_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14586_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14586_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11798_ _11798_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__or2_1
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ _13537_/A _13537_/B vssd1 vssd1 vccd1 vccd1 _15597_/D sky130_fd_sc_hd__xor2_1
X_10749_ _15716_/Q _15782_/Q vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__or2_1
XFILLER_9_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12953__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater535_A _13826_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _13468_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _13470_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__15686__D _15686_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15207_ _15367_/CLK _15207_/D _14254_/Y vssd1 vssd1 vccd1 vccd1 _15207_/Q sky130_fd_sc_hd__dfrtp_1
X_12419_ _12420_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater702_A _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07579__A0 _15475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13399_ _13399_/A _13411_/A vssd1 vssd1 vccd1 vccd1 _13400_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _15400_/CLK _15138_/D _14181_/Y vssd1 vssd1 vccd1 vccd1 _15138_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07960_ _07960_/A _10963_/A vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__nor2_1
X_15069_ _15345_/CLK _15069_/D _14108_/Y vssd1 vssd1 vccd1 vccd1 _15069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15571_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08878__A _15468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07891_ _07891_/A vssd1 vssd1 vccd1 vccd1 _15322_/D sky130_fd_sc_hd__clkbuf_1
X_09630_ _09630_/A vssd1 vssd1 vccd1 vccd1 _15301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _09783_/A _09561_/B vssd1 vssd1 vccd1 vccd1 _15173_/D sky130_fd_sc_hd__xor2_1
XFILLER_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08512_ _14917_/Q vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__buf_4
XFILLER_70_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _09535_/A _09492_/B vssd1 vssd1 vccd1 vccd1 _15282_/D sky130_fd_sc_hd__xnor2_1
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08466_/C sky130_fd_sc_hd__xor2_1
XFILLER_93_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08374_ _08728_/B _12627_/A _08391_/A _08373_/X vssd1 vssd1 vccd1 vccd1 _08404_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08118__A _08118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07806__A1 input169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13959__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11479__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_896 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__B _15029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13107__A2 _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09828_ _15057_/Q _09827_/Y _09826_/B vssd1 vssd1 vccd1 vccd1 _09830_/B sky130_fd_sc_hd__a21o_1
XFILLER_48_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08298__A1 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A x_i_7[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _08702_/A _13636_/A _12769_/A _13645_/B _12625_/X vssd1 vssd1 vccd1 vccd1
+ _12771_/B sky130_fd_sc_hd__a221o_1
XANTENNA__08298__B2 _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12381_/A _11721_/B vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__xnor2_4
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__buf_6
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11652_ _12372_/B _11652_/B vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__xor2_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08028__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10603_ _10527_/A _10602_/B _10527_/B vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__a21boi_1
XFILLER_156_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _14376_/A vssd1 vssd1 vccd1 vccd1 _14371_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__or2_1
XFILLER_210_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13322_ _13491_/S _13322_/B vssd1 vssd1 vccd1 vccd1 _13325_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input81_A x_i_4[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10534_ _10532_/Y _10534_/B vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__and2b_1
XFILLER_122_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09067__B_N _15478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__A _15757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ _15127_/Q _10464_/Y _10463_/B vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__a21o_1
X_13253_ _13422_/A _13253_/B vssd1 vssd1 vccd1 vccd1 _13300_/A sky130_fd_sc_hd__and2_1
XFILLER_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__or2_1
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ _10395_/B _10395_/C _10395_/A vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__o21ai_1
X_13184_ _13366_/A vssd1 vssd1 vccd1 vccd1 _13253_/B sky130_fd_sc_hd__inv_2
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12244_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__or2_1
XFILLER_2_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07806__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11836__B _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _12312_/S _12247_/A _12244_/A vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__and3_1
XFILLER_172_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output335_A _11352_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater708 _07536_/S vssd1 vssd1 vccd1 vccd1 _07538_/S sky130_fd_sc_hd__buf_6
Xrepeater719 _15700_/Q vssd1 vssd1 vccd1 vccd1 output394/A sky130_fd_sc_hd__clkbuf_2
X_11017_ _14988_/Q _14922_/Q vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13109__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ _15758_/CLK _15756_/D _14834_/Y vssd1 vssd1 vccd1 vccd1 _15756_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12968_ _12867_/A _12966_/X _12967_/X vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__a21oi_2
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14707_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _11920_/A _11920_/B vssd1 vssd1 vccd1 vccd1 _11921_/A sky130_fd_sc_hd__or2_1
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15687_ _15687_/CLK _15687_/D _14761_/Y vssd1 vssd1 vccd1 vccd1 _15687_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ _12940_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__xnor2_1
XFILLER_127_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14638_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09789__A1 _15436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14569_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14569_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater917_A input193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__nand2_1
XFILLER_140_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15666__CLK _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08992_ _13597_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _15105_/D sky130_fd_sc_hd__xor2_1
XANTENNA__14403__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _15119_/Q _15152_/Q vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__or2_1
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07874_ _15330_/Q input135/X _07892_/S vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _09613_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _15181_/D sky130_fd_sc_hd__nor2_1
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12858__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09544_ _15431_/Q _15415_/Q vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07451__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09475_ _09473_/X _09480_/B vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__and2b_1
XFILLER_169_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10378__A _15135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08426_ _08426_/A _08426_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ _12810_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08369_/A sky130_fd_sc_hd__nand2_1
XFILLER_211_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08790__B _15323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08288_ _08288_/A _08288_/B vssd1 vssd1 vccd1 vccd1 _08289_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10250_ _15079_/Q _15244_/Q vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__or2b_1
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11937__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _15315_/Q _15150_/Q vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__and2b_1
XFILLER_191_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14313__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07626__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13940_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13940_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input233_A x_r_6[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13871_ _14985_/Q _13871_/B vssd1 vssd1 vccd1 vccd1 _13871_/X sky130_fd_sc_hd__or2_1
XFILLER_19_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15610_ _15705_/CLK _15610_/D _14680_/Y vssd1 vssd1 vccd1 vccd1 _15610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12822_ _12921_/A _12881_/A vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09142__A _15562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15572_/CLK _15541_/D _14607_/Y vssd1 vssd1 vccd1 vccd1 _15541_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _12799_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _12779_/A sky130_fd_sc_hd__xnor2_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11733_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15472_/CLK _15472_/D _14534_/Y vssd1 vssd1 vccd1 vccd1 _15472_/Q sky130_fd_sc_hd__dfrtp_1
X_12684_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__or2_1
XFILLER_70_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_525 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14423_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14423_/Y sky130_fd_sc_hd__inv_2
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14354_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14354_/Y sky130_fd_sc_hd__inv_2
X_11566_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__xor2_1
XFILLER_183_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output285_A output285/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _13350_/A _13305_/B vssd1 vssd1 vccd1 vccd1 _13307_/A sky130_fd_sc_hd__xnor2_1
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10517_ _15255_/Q _10516_/Y _10512_/B vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14285_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14285_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12008__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _12360_/B _11507_/B vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__xnor2_4
XFILLER_196_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13236_ _13157_/A _13157_/B _13235_/X vssd1 vssd1 vccd1 vccd1 _13238_/B sky130_fd_sc_hd__a21o_1
XFILLER_170_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10448_ _15156_/Q vssd1 vssd1 vccd1 vccd1 _10448_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output452_A output452/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13219_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14223__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ _10379_/A _10486_/A vssd1 vssd1 vccd1 vccd1 _15791_/D sky130_fd_sc_hd__xnor2_1
XFILLER_124_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07536__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12118_ _12119_/A _12119_/B _12119_/C vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09317__A _15391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13098_ _13098_/A _13206_/A vssd1 vssd1 vccd1 vccd1 _13100_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _12050_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _12119_/B sky130_fd_sc_hd__and2_1
Xrepeater538 _11298_/X vssd1 vssd1 vccd1 vccd1 output470/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater549 repeater550/X vssd1 vssd1 vccd1 vccd1 output467/A sky130_fd_sc_hd__buf_6
XANTENNA_repeater867_A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__B _15450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15808_ _15808_/CLK _15808_/D _14888_/Y vssd1 vssd1 vccd1 vccd1 _15808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07590_ _07590_/A vssd1 vssd1 vccd1 vccd1 _15470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_959 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15739_ _15741_/CLK _15739_/D _14816_/Y vssd1 vssd1 vccd1 vccd1 _15739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _15246_/D sky130_fd_sc_hd__nor2_1
XFILLER_178_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08211_/X sky130_fd_sc_hd__or2_1
XFILLER_53_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09191_ _09191_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _15294_/D sky130_fd_sc_hd__nor2_1
XFILLER_178_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13302__A _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ _15016_/Q vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__buf_6
XFILLER_193_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08073_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11806_/C sky130_fd_sc_hd__inv_2
XFILLER_105_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14133__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08975_ _15475_/Q _15459_/Q _08974_/X vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13972__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07926_ _15053_/Q _15086_/Q vssd1 vssd1 vccd1 vccd1 _07927_/B sky130_fd_sc_hd__or2_1
XFILLER_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07857_ _07857_/A vssd1 vssd1 vccd1 vccd1 _15339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09237__A_N _15499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07788_ _07788_/A vssd1 vssd1 vccd1 vccd1 _15373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ _15537_/Q _15521_/Q vssd1 vssd1 vccd1 vccd1 _09527_/X sky130_fd_sc_hd__and2_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09458_/A _09466_/A vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08391_/A _08391_/B _08408_/X vssd1 vssd1 vccd1 vccd1 _08432_/A sky130_fd_sc_hd__o21ai_1
XFILLER_12_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14953__D _14953_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09389_ _09389_/A vssd1 vssd1 vccd1 vccd1 _15146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14308__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11420_ _11418_/A _11418_/B _11419_/X vssd1 vssd1 vccd1 vccd1 _11421_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10232__A1 _15075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _11350_/A _11350_/B _11099_/B vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__a21oi_2
XANTENNA_input183_A x_r_3[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _15122_/Q _15155_/Q vssd1 vssd1 vccd1 vccd1 _10304_/A sky130_fd_sc_hd__or2_1
X_14070_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14070_/Y sky130_fd_sc_hd__inv_2
X_11282_ _15784_/Q _15718_/Q vssd1 vssd1 vccd1 vccd1 _11283_/C sky130_fd_sc_hd__or2b_1
XANTENNA__15784__D _15784_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11667__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13021_ _13021_/A _13021_/B vssd1 vssd1 vccd1 vccd1 _13022_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10233_ _11404_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _15765_/D sky130_fd_sc_hd__xor2_1
XFILLER_156_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14043__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _15147_/Q _15312_/Q vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input44_A x_i_2[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__B _15034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14972_ _15508_/CLK _14972_/D _14005_/Y vssd1 vssd1 vccd1 vccd1 _14972_/Q sky130_fd_sc_hd__dfrtp_1
X_10095_ _15216_/Q _15117_/Q vssd1 vssd1 vccd1 vccd1 _10095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13923_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13849_/X _13850_/X _13851_/X _13853_/X _13767_/B vssd1 vssd1 vccd1 vccd1
+ _13859_/B sky130_fd_sc_hd__o41a_1
XFILLER_63_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12805_ _12805_/A _12805_/B _12805_/C vssd1 vssd1 vccd1 vccd1 _13056_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13106__B _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13785_ _13785_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13867_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10997_ _10997_/A vssd1 vssd1 vccd1 vccd1 _15013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15524_ _15561_/CLK _15524_/D _14589_/Y vssd1 vssd1 vccd1 vccd1 _15524_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12736_ _12670_/A _12670_/B _12735_/X vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__a21bo_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15455_ _15573_/CLK _15455_/D _14516_/Y vssd1 vssd1 vccd1 vccd1 _15455_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _13046_/A _12871_/A _12667_/C vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__and3_1
XANTENNA__14218__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__inv_2
X_11618_ _11561_/B _11618_/B vssd1 vssd1 vccd1 vccd1 _11618_/X sky130_fd_sc_hd__and2b_1
XFILLER_129_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15386_ _15808_/CLK _15386_/D _14444_/Y vssd1 vssd1 vccd1 vccd1 _15386_/Q sky130_fd_sc_hd__dfrtp_1
X_12598_ _12596_/A _12433_/B _12596_/B _12431_/X vssd1 vssd1 vccd1 vccd1 _12599_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14337_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14337_/Y sky130_fd_sc_hd__inv_2
X_11549_ _11620_/B _11549_/B vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__xnor2_1
XFILLER_183_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14268_ _14269_/A vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15694__D _15694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13219_ _13219_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__or2b_1
XFILLER_48_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14199_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14218_/A sky130_fd_sc_hd__buf_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14888__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_clk clkbuf_1_1_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08760_ _15318_/Q _15334_/Q vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__and2b_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07711_ _07711_/A vssd1 vssd1 vccd1 vccd1 _15411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08691_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _08692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_211_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11516__S _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07642_ _15444_/Q _07642_/A1 _07644_/S vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07573_ _15478_/Q _07573_/A1 _07591_/S vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _15406_/Q _15390_/Q vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__and2_1
XFILLER_94_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09243_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__and2_1
XANTENNA__10656__A _15273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14128__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _15567_/Q _15547_/Q _09173_/X vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__a21oi_1
XFILLER_182_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _15009_/Q vssd1 vssd1 vccd1 vccd1 _11707_/A sky130_fd_sc_hd__buf_6
XFILLER_175_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13967__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__A _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11962__A1 _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08056_ _11435_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08057_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13686__B _13824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12911__B1 _12910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14798__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput105 x_i_6[15] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07394__A1 input130/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 x_i_7[10] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput127 x_i_7[6] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13467__A1 _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08958_ _08890_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _08959_/C sky130_fd_sc_hd__and2b_1
Xinput138 x_r_0[1] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput149 x_r_1[11] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__clkbuf_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ _07909_/A vssd1 vssd1 vccd1 vccd1 _15185_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14948__D _14948_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _15470_/Q _15454_/Q vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__and2_1
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _14897_/Q _14963_/Q vssd1 vssd1 vccd1 vccd1 _10924_/B sky130_fd_sc_hd__or2b_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater880 input247/X vssd1 vssd1 vccd1 vccd1 _07647_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater891 input233/X vssd1 vssd1 vccd1 vccd1 _07773_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10851_ _10850_/A _10850_/B _10167_/B vssd1 vssd1 vccd1 vccd1 _10852_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13570_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _13571_/B sky130_fd_sc_hd__nor2_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/A vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15779__D _15779_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ _12332_/A _12332_/B _12520_/Y vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__a21o_1
XFILLER_9_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14038__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15240_ _15347_/CLK _15240_/D _14289_/Y vssd1 vssd1 vccd1 vccd1 _15240_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12440_/A _12455_/C _12451_/X vssd1 vssd1 vccd1 vccd1 _12456_/B sky130_fd_sc_hd__a21oi_1
XFILLER_200_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11403_ _10221_/Y _11402_/B _10223_/B vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__08949__A2 _15450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15171_ _15433_/CLK _15171_/D _14215_/Y vssd1 vssd1 vccd1 vccd1 _15171_/Q sky130_fd_sc_hd__dfrtp_1
X_12383_ _12391_/C _12389_/C _12384_/A vssd1 vssd1 vccd1 vccd1 _12383_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14122_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14122_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11334_ _14996_/Q _14930_/Q vssd1 vssd1 vccd1 vccd1 _11335_/C sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_55_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14053_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14053_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11265_ _11265_/A _11265_/B vssd1 vssd1 vccd1 vccd1 _11267_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13004_ _13072_/A _13071_/A vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10216_ _10216_/A _10216_/B vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__nand2_2
X_11196_ _11195_/A _11195_/C _11367_/A vssd1 vssd1 vccd1 vccd1 _11197_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__15019__D _15019_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10147_ _10147_/A _10843_/A vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13458__A1 _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07814__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_113_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1062 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14955_ _15184_/CLK _14955_/D _13987_/Y vssd1 vssd1 vccd1 vccd1 _14955_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__nor2_2
XANTENNA_output415_A output415/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _15345_/Q _15329_/Q vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and2_1
X_14886_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14886_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13837_ _13837_/A vssd1 vssd1 vccd1 vccd1 _13838_/A sky130_fd_sc_hd__inv_2
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_128_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13768_ _14983_/Q vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__inv_2
XFILLER_189_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12675__B _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12719_ _12643_/A _12643_/B _12718_/Y vssd1 vssd1 vccd1 vccd1 _12811_/B sky130_fd_sc_hd__a21o_1
X_15507_ _15572_/CLK _15507_/D _14571_/Y vssd1 vssd1 vccd1 vccd1 _15507_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_repeater732_A repeater733/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_13699_ _13696_/A _13826_/A _13698_/X vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__a21o_1
XFILLER_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15438_ _15438_/CLK _15438_/D _14498_/Y vssd1 vssd1 vccd1 vccd1 _15438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15749_/CLK _15369_/D _14425_/Y vssd1 vssd1 vccd1 vccd1 _15369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _15228_/Q _15195_/Q vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__or2b_1
XFILLER_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _15756_/D sky130_fd_sc_hd__xor2_1
XFILLER_140_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08811_/A _08811_/B _13897_/B vssd1 vssd1 vccd1 vccd1 _08818_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09572_/Y _09791_/B _09574_/B vssd1 vssd1 vccd1 vccd1 _09794_/B sky130_fd_sc_hd__o21ai_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14411__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07724__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08739_/X _08740_/X _08741_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _08743_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13027__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09224__B _09224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _12688_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08675_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07625_ _07625_/A vssd1 vssd1 vccd1 vccd1 _15453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07556_ _07556_/A vssd1 vssd1 vccd1 vccd1 _15487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13621__A1 _15376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15599__D _15599_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _07699_/A vssd1 vssd1 vccd1 vccd1 _07536_/S sky130_fd_sc_hd__buf_8
XFILLER_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09226_ _09225_/Y _15479_/Q _09224_/B vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__a21o_1
XFILLER_167_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _09636_/A _09157_/B vssd1 vssd1 vccd1 vccd1 _15287_/D sky130_fd_sc_hd__xor2_1
X_08108_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _09086_/Y _09088_/B vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__nand2b_2
XFILLER_123_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08039_ _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__xor2_1
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_502 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09575__A_N _15436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11050_ _11042_/Y _11046_/B _11044_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__o21ai_2
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ _15198_/Q _15231_/Q vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__and2_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14321__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input146_A x_r_0[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09108__A2 _15485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14740_/Y sky130_fd_sc_hd__inv_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11952_ _12426_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _11952_/Y sky130_fd_sc_hd__nand2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09134__B _15492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10903_ _10902_/A _10902_/C _11117_/A vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__o21ai_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14671_/Y sky130_fd_sc_hd__inv_2
X_11883_ _12055_/A _11977_/A _11898_/A vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__and3b_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13622_ _13622_/A _13622_/B vssd1 vssd1 vccd1 vccd1 _15098_/D sky130_fd_sc_hd__xor2_1
X_10834_ _10834_/A _10834_/B _10834_/C vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__or3_1
XFILLER_38_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09150__A _15563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _15764_/Q vssd1 vssd1 vccd1 vccd1 _13553_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10296__A _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ _15785_/Q _15719_/Q vssd1 vssd1 vccd1 vccd1 _11287_/A sky130_fd_sc_hd__or2b_1
XFILLER_185_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12504_ _14951_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12504_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13484_ _13781_/B _13781_/A vssd1 vssd1 vccd1 vccd1 _13484_/X sky130_fd_sc_hd__and2b_1
X_10696_ _15181_/Q _15280_/Q vssd1 vssd1 vccd1 vccd1 _10697_/B sky130_fd_sc_hd__and2b_1
XFILLER_157_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15223_ _15498_/CLK _15223_/D _14271_/Y vssd1 vssd1 vccd1 vccd1 _15223_/Q sky130_fd_sc_hd__dfrtp_1
X_12435_ _12435_/A _12435_/B _12597_/A vssd1 vssd1 vccd1 vccd1 _12436_/B sky130_fd_sc_hd__or3b_1
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15154_ _15279_/CLK _15154_/D _14197_/Y vssd1 vssd1 vccd1 vccd1 _15154_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11839__B _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _12366_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__nor2_1
Xoutput409 output409/A vssd1 vssd1 vccd1 vccd1 y_r_0[6] sky130_fd_sc_hd__buf_2
XANTENNA_output365_A output365/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14105_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15085_ _15347_/CLK _15085_/D _14125_/Y vssd1 vssd1 vccd1 vccd1 _15085_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12297_ _15739_/Q _12304_/B vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__nor2_1
X_14036_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__inv_2
X_11248_ _11248_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _11248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14231__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _11177_/Y _11179_/B vssd1 vssd1 vccd1 vccd1 _11363_/A sky130_fd_sc_hd__and2b_2
XFILLER_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater682_A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14938_ _15464_/CLK _14938_/D _13969_/Y vssd1 vssd1 vccd1 vccd1 _14938_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_208_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14869_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14869_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07530__A1 input111/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _15562_/Q _07410_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__mux2_1
X_08390_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ _13605_/A _09008_/B _09010_/X vssd1 vssd1 vccd1 vccd1 _09012_/B sky130_fd_sc_hd__a21o_1
XFILLER_192_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10934__A _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14406__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09913_ _09983_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09844_ _15061_/Q _09843_/Y _09842_/B vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__a21o_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14141__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09775_ _09775_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _15154_/D sky130_fd_sc_hd__xnor2_1
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_550 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13980__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1060 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08726_ _12810_/A _12780_/A vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__xnor2_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__xor2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _15461_/Q input67/X _07632_/S vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08588_ _08711_/B vssd1 vssd1 vccd1 vccd1 _08588_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07539_ _07539_/A vssd1 vssd1 vccd1 vccd1 _15495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ _10550_/A _10558_/A vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__nand2_1
XFILLER_195_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _15576_/Q _15556_/Q vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__and2_1
XFILLER_185_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14961__D _14961_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10481_ _10480_/A _10480_/B _10359_/B vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__a21o_1
XFILLER_154_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14316__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ _12220_/A _12220_/B vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__or2_1
XFILLER_136_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13220__A _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12151_ _12466_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12456_/A sky130_fd_sc_hd__xor2_1
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11102_ _11100_/A _11350_/A _11101_/Y vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__and2_1
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11033_ _14925_/Q _14991_/Q vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14051__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12884__A2 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _12985_/C _12985_/B _13020_/B vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__a21boi_1
X_15772_ _15773_/CLK _15772_/D _14851_/Y vssd1 vssd1 vccd1 vccd1 _15772_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11935_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__nand2_1
X_14723_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14723_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07512__A1 _07512_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14654_/Y sky130_fd_sc_hd__inv_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11866_/A _11866_/B _11866_/C _11866_/D vssd1 vssd1 vccd1 vccd1 _11867_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_33_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13605_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _15092_/D sky130_fd_sc_hd__xor2_1
XFILLER_32_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10817_ _10817_/A _10817_/B vssd1 vssd1 vccd1 vccd1 _14908_/D sky130_fd_sc_hd__xor2_1
XFILLER_207_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14585_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14585_/Y sky130_fd_sc_hd__inv_2
X_11797_ _11797_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13536_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13537_/B sky130_fd_sc_hd__and2_1
XFILLER_186_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10748_ _11267_/A _10748_/B vssd1 vssd1 vccd1 vccd1 _10748_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output482_A output482/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12953__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ _13352_/A _13417_/B _13354_/B vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__o21a_1
XFILLER_199_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10679_ _10679_/A _10679_/B vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__nand2_2
XANTENNA__14226__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15206_ _15367_/CLK _15206_/D _14253_/Y vssd1 vssd1 vccd1 vccd1 _15206_/Q sky130_fd_sc_hd__dfrtp_1
X_12418_ _12418_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13398_ _13399_/A _13411_/A vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__or2_1
XFILLER_154_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07579__A1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15137_ _15400_/CLK _15137_/D _14180_/Y vssd1 vssd1 vccd1 vccd1 _15137_/Q sky130_fd_sc_hd__dfrtp_1
X_12349_ _12332_/A _12331_/A _12348_/X vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__o21a_1
XFILLER_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15068_ _15346_/CLK _15068_/D _14107_/Y vssd1 vssd1 vccd1 vccd1 _15068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater897_A repeater898/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__B _15452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14019_/Y sky130_fd_sc_hd__inv_2
X_07890_ _15322_/Q _07890_/A1 _07892_/S vssd1 vssd1 vccd1 vccd1 _07891_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15207__D _15207_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09560_ _09781_/A _09557_/B _09559_/X vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _13390_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_695 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09491_ _09490_/Y _15523_/Q _09486_/B vssd1 vssd1 vccd1 vccd1 _09492_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _08462_/A _08462_/B _08464_/A vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__or3_1
XFILLER_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _12810_/A _08369_/B _08421_/B vssd1 vssd1 vccd1 vccd1 _08373_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14136__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13975__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09827_ _15090_/Q vssd1 vssd1 vccd1 vccd1 _09827_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07742__A1 _07742_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _15100_/Q _15067_/Q vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__and2b_1
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11241__B_N _15757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08709_ _08713_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__nand2_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11942__B _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08298__A2 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _15054_/Q _15087_/Q _09687_/Y _09688_/Y vssd1 vssd1 vccd1 vccd1 _09693_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ _11651_/A _11651_/B _11718_/X _11719_/X vssd1 vssd1 vccd1 vccd1 _11721_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input109_A x_i_6[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11651_ _11651_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__nand2_1
XFILLER_199_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10602_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _14994_/D sky130_fd_sc_hd__xnor2_1
XFILLER_168_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14370_ _14376_/A vssd1 vssd1 vccd1 vccd1 _14370_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _11580_/A _12529_/A _11581_/X vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__a21o_1
XFILLER_156_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ _13321_/A vssd1 vssd1 vccd1 vccd1 _13322_/B sky130_fd_sc_hd__inv_2
XFILLER_127_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ _15259_/Q _15292_/Q vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_734 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14046__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_907 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ _13253_/B _13357_/B _13273_/A vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__and3_1
XFILLER_202_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10464_ _15160_/Q vssd1 vssd1 vccd1 vccd1 _10464_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input74_A x_i_4[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11389__B _15035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13183_/A _13273_/A _13201_/A vssd1 vssd1 vccd1 vccd1 _13187_/A sky130_fd_sc_hd__and3_1
XFILLER_89_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10395_ _10395_/A _10395_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__or3_1
XFILLER_159_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12134_ _12244_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12065_ _12312_/S _12244_/A _12247_/A vssd1 vssd1 vccd1 vccd1 _12075_/A sky130_fd_sc_hd__a21oi_1
XFILLER_123_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater709 _07536_/S vssd1 vssd1 vccd1 vccd1 _07532_/S sky130_fd_sc_hd__buf_4
X_11016_ _11016_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _15020_/D sky130_fd_sc_hd__xnor2_1
XFILLER_65_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output328_A output328/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07822__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _12967_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12967_/X sky130_fd_sc_hd__and2_1
X_15755_ _15758_/CLK _15755_/D _14833_/Y vssd1 vssd1 vccd1 vccd1 _15755_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11918_ _11986_/A _11985_/A vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__xor2_1
X_14706_ _14709_/A vssd1 vssd1 vccd1 vccd1 _14706_/Y sky130_fd_sc_hd__inv_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15686_ _15687_/CLK _15686_/D _14760_/Y vssd1 vssd1 vccd1 vccd1 _15686_/Q sky130_fd_sc_hd__dfrtp_1
X_12898_ _12826_/A _12826_/B _12820_/A vssd1 vssd1 vccd1 vccd1 _12940_/B sky130_fd_sc_hd__a21o_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _11928_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__nand2_1
X_14637_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14637_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater645_A _10723_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09789__A2 _15420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14568_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14568_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater812_A _15577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ _13803_/A _13519_/B vssd1 vssd1 vccd1 vccd1 _13519_/Y sky130_fd_sc_hd__nand2_1
X_14499_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14499_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13795__A _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08889__A _15470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12821__B1_N _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_718 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08991_ _08990_/Y _15351_/Q _08988_/B vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _15119_/Q _15152_/Q vssd1 vssd1 vccd1 vccd1 _10295_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12204__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _07873_/A vssd1 vssd1 vccd1 vccd1 _15331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_818 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07724__A1 input224/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09612_ _09611_/A _09611_/B _09806_/A vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07732__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09543_ _09545_/B _09543_/B vssd1 vssd1 vccd1 vccd1 _15169_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09474_ _09473_/A _09473_/B _09526_/A vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08129__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08425_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08426_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09016__A_N _15372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ _15037_/Q vssd1 vssd1 vccd1 vccd1 _12627_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_149_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08287_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08287_/X sky130_fd_sc_hd__xor2_1
XFILLER_177_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07412__A0 _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _15150_/Q _15315_/Q vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__and2b_1
XFILLER_161_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11511__A2 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _14985_/Q _13871_/B vssd1 vssd1 vccd1 vccd1 _13870_/X sky130_fd_sc_hd__and2_1
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input226_A x_r_5[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07642__S _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ _13201_/A _12714_/B _13012_/A vssd1 vssd1 vccd1 vccd1 _12825_/A sky130_fd_sc_hd__a21boi_1
XFILLER_75_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12800_/A _12800_/B vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__xnor2_1
X_15540_ _15573_/CLK _15540_/D _14606_/Y vssd1 vssd1 vccd1 vccd1 _15540_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11634_/A _11633_/B _11633_/A vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__o21bai_1
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15471_ _15558_/CLK _15471_/D _14533_/Y vssd1 vssd1 vccd1 vccd1 _15471_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12683_/A _12683_/B vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__xnor2_1
XFILLER_188_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14422_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14422_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11634_ _11634_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14353_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14353_/Y sky130_fd_sc_hd__inv_2
X_11565_ _11563_/Y _11487_/B _11564_/X vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__o21a_1
XFILLER_129_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13304_ _13356_/A _13350_/C vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__nor2_1
X_10516_ _15288_/Q vssd1 vssd1 vccd1 vccd1 _10516_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14284_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14284_/Y sky130_fd_sc_hd__inv_2
X_11496_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11507_/B sky130_fd_sc_hd__xnor2_4
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output278_A output278/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _13156_/B _13235_/B vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__and2b_1
XFILLER_196_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10447_ _10447_/A _10447_/B vssd1 vssd1 vccd1 vccd1 _14892_/D sky130_fd_sc_hd__nor2_1
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14504__A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13166_ _13118_/A _13118_/B _13165_/X vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__o21ai_1
X_10378_ _15135_/Q _15168_/Q vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__xnor2_2
XFILLER_123_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output445_A output445/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12117_ _12117_/A _12161_/A vssd1 vssd1 vccd1 vccd1 _12119_/C sky130_fd_sc_hd__xnor2_1
XFILLER_170_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13097_ _13097_/A _13097_/B _13097_/C vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__nand3_1
XFILLER_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12048_ _11966_/A _11966_/B _11963_/X vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__a21o_1
XFILLER_133_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07706__A1 _07706_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater595_A _11321_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater539 _11243_/Y vssd1 vssd1 vccd1 vccd1 output504/A sky130_fd_sc_hd__buf_4
XFILLER_172_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15807_ _15808_/CLK _15807_/D _14887_/Y vssd1 vssd1 vccd1 vccd1 _15807_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ _14003_/A vssd1 vssd1 vccd1 vccd1 _13999_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15738_ _15790_/CLK _15738_/D _14815_/Y vssd1 vssd1 vccd1 vccd1 _15738_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ _15771_/CLK _15669_/D _14743_/Y vssd1 vssd1 vccd1 vccd1 _15669_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__xnor2_1
XFILLER_194_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07890__A0 _15322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09190_ _09189_/A _09189_/C _09659_/A vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__o21a_1
XFILLER_147_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08141_ _08139_/A _08236_/B _08140_/X vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__a21bo_1
XFILLER_147_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ _15801_/Q vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__buf_4
XFILLER_101_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14414__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08974_ _15475_/Q _15459_/Q _08973_/B vssd1 vssd1 vccd1 vccd1 _08974_/X sky130_fd_sc_hd__o21a_1
XFILLER_29_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07925_ _15053_/Q _15086_/Q vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nand2_1
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07856_ _15339_/Q input207/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07857_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _15373_/Q input241/X _07791_/S vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09526_ _09526_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _15263_/D sky130_fd_sc_hd__xor2_1
XFILLER_71_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09457_ _15535_/Q _15519_/Q vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__or2b_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09870__A1 _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08408_/X sky130_fd_sc_hd__or2_1
XFILLER_196_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09388_ _09386_/X _09390_/C vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__and2b_1
XFILLER_178_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08339_ _08327_/X _08285_/Y _08328_/Y _08289_/X _08338_/X vssd1 vssd1 vccd1 vccd1
+ _08339_/X sky130_fd_sc_hd__a221o_1
XFILLER_184_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12109__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15130__D _15130_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11091__A_N _15001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _11350_/A _11350_/B vssd1 vssd1 vccd1 vccd1 _11350_/X sky130_fd_sc_hd__xor2_1
XFILLER_137_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ _10301_/A _10437_/B vssd1 vssd1 vccd1 vccd1 _15777_/D sky130_fd_sc_hd__xnor2_1
XFILLER_192_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11281_ _11281_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14324__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input176_A x_r_2[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _13020_/A _13020_/B vssd1 vssd1 vccd1 vccd1 _13022_/C sky130_fd_sc_hd__nor2_1
XFILLER_152_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10232_ _15075_/Q _10231_/Y _10227_/B vssd1 vssd1 vccd1 vccd1 _10234_/B sky130_fd_sc_hd__a21o_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ _10163_/A vssd1 vssd1 vccd1 vccd1 _15804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input37_A x_i_2[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _15508_/CLK _14971_/D _14004_/Y vssd1 vssd1 vccd1 vccd1 _14971_/Q sky130_fd_sc_hd__dfrtp_1
X_10094_ _10094_/A _10432_/A vssd1 vssd1 vccd1 vccd1 _14985_/D sky130_fd_sc_hd__xor2_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13922_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13922_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_607 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13853_ _13752_/A _13752_/B _13842_/C _13852_/Y _13842_/A vssd1 vssd1 vccd1 vccd1
+ _13853_/X sky130_fd_sc_hd__o221a_1
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12804_ _12805_/A _12805_/B _12805_/C vssd1 vssd1 vccd1 vccd1 _12804_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ _10996_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__and2_1
X_13784_ _13772_/B _13772_/C _13783_/X _13771_/B vssd1 vssd1 vccd1 vccd1 _13785_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12996__A1 _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15523_ _15528_/CLK _15523_/D _14588_/Y vssd1 vssd1 vccd1 vccd1 _15523_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12803_/A _12735_/B _12735_/C vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__or3_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07872__A0 _15331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15454_ _15727_/CLK _15454_/D _14515_/Y vssd1 vssd1 vccd1 vccd1 _15454_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12803_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__nor2_1
XFILLER_203_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output395_A output395/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14405_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14405_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12597_ _12597_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _15684_/D sky130_fd_sc_hd__xnor2_1
X_15385_ _15803_/CLK _15385_/D _14443_/Y vssd1 vssd1 vccd1 vccd1 _15385_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__15040__D _15040_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ _11622_/A _08144_/A _11707_/A vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__mux2_1
X_14336_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14336_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14267_ _14269_/A vssd1 vssd1 vccd1 vccd1 _14267_/Y sky130_fd_sc_hd__inv_2
X_11479_ _11707_/A _11746_/A vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater608_A _11264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14234__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ _13210_/A _13715_/A _13217_/Y vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07547__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _13491_/S _14920_/Q vssd1 vssd1 vccd1 vccd1 _13150_/C sky130_fd_sc_hd__nor2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater977_A input115/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ _15411_/Q input216/X _07750_/S vssd1 vssd1 vccd1 vccd1 _07711_/A sky130_fd_sc_hd__mux2_1
X_08690_ _08526_/A _08526_/B _08689_/Y vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07641_ _07641_/A vssd1 vssd1 vccd1 vccd1 _15445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11239__A1 _15756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ _07572_/A vssd1 vssd1 vccd1 vccd1 _15479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09311_ _15406_/Q _15390_/Q vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14409__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _15242_/D sky130_fd_sc_hd__xor2_2
XFILLER_178_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09173_ _15567_/Q _15547_/Q _09169_/B vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__o21a_1
X_08124_ _15005_/Q vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__buf_4
XFILLER_193_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_929 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ _08058_/A _08058_/B vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__xor2_2
XFILLER_135_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14144__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07457__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13983__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 x_i_6[1] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07981__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput117 x_i_7[11] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_1
Xinput128 x_i_7[7] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_2
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput139 x_r_0[2] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _08957_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _15194_/D sky130_fd_sc_hd__xnor2_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07908_ _08936_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__and2_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _15470_/Q _15454_/Q vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__nor2_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater870 input32/X vssd1 vssd1 vccd1 vccd1 _07496_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07839_ _07839_/A vssd1 vssd1 vccd1 vccd1 _15348_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater881 input245/X vssd1 vssd1 vccd1 vccd1 _07651_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater892 input231/X vssd1 vssd1 vccd1 vccd1 _07777_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10850_ _10850_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _14917_/D sky130_fd_sc_hd__xor2_2
XFILLER_186_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11950__B _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09509_/A _09509_/B vssd1 vssd1 vccd1 vccd1 _15257_/D sky130_fd_sc_hd__xor2_1
X_10781_ _10779_/X _10787_/A vssd1 vssd1 vccd1 vccd1 _10781_/X sky130_fd_sc_hd__and2b_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14319__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _12520_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12520_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13223__A _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ _12105_/B _12451_/B vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__and2b_1
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07606__A0 _15462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _15732_/D sky130_fd_sc_hd__xnor2_2
X_15170_ _15170_/CLK _15170_/D _14214_/Y vssd1 vssd1 vccd1 vccd1 _15170_/Q sky130_fd_sc_hd__dfrtp_1
X_12382_ _14942_/Q vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__inv_2
XFILLER_197_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15795__D _15795_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11678__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _11333_/A _11333_/B vssd1 vssd1 vccd1 vccd1 _11335_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14054__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14052_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _11265_/A _11265_/B vssd1 vssd1 vccd1 vccd1 _11264_/X sky130_fd_sc_hd__xor2_4
XFILLER_141_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13003_ _13086_/A _13086_/B vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10215_ _15074_/Q _15239_/Q vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11195_ _11195_/A _11367_/A _11195_/C vssd1 vssd1 vccd1 vccd1 _11197_/A sky130_fd_sc_hd__and3_1
XFILLER_80_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _15310_/Q _15145_/Q vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__or2b_1
XFILLER_39_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14954_ _15791_/CLK _14954_/D _13986_/Y vssd1 vssd1 vccd1 vccd1 _14954_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10077_ _15115_/Q _15214_/Q vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__and2b_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08334__A1 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13905_ _13905_/A _13905_/B vssd1 vssd1 vccd1 vccd1 _15065_/D sky130_fd_sc_hd__xor2_1
XANTENNA_output310_A _10918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14885_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output408_A output408/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ _13836_/A _13836_/B vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__or2_1
XFILLER_46_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07830__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_662 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10979_ _10980_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _15009_/D sky130_fd_sc_hd__xor2_1
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _15704_/D sky130_fd_sc_hd__xor2_1
XFILLER_206_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14229__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater558_A _11137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15506_/CLK _15506_/D _14570_/Y vssd1 vssd1 vccd1 vccd1 _15506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12718_ _12718_/A _12718_/B vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_203_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13698_ _13827_/B _14976_/Q vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__and2b_1
X_15437_ _15437_/CLK _15437_/D _14497_/Y vssd1 vssd1 vccd1 vccd1 _15437_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12649_ _12726_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_851 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15368_ _15374_/CLK _15368_/D _14424_/Y vssd1 vssd1 vccd1 vccd1 _15368_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14319_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15299_ _15572_/CLK _15299_/D _14351_/Y vssd1 vssd1 vccd1 vccd1 _15299_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09860_ _09859_/A _09859_/B _09751_/B vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__a21o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08897__A _15455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _08811_/A _08811_/B _13897_/B vssd1 vssd1 vccd1 vccd1 _08811_/X sky130_fd_sc_hd__and3_1
XFILLER_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09791_ _09791_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _15160_/D sky130_fd_sc_hd__xor2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08601_/X _08742_/B vssd1 vssd1 vccd1 vccd1 _08742_/X sky130_fd_sc_hd__and2b_1
XFILLER_100_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12212__A _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13027__B _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ _08524_/A _08539_/B _08672_/X vssd1 vssd1 vccd1 vccd1 _08692_/A sky130_fd_sc_hd__a21bo_1
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07624_ _15453_/Q _07624_/A1 _07644_/S vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07740__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07555_ _15487_/Q _07555_/A1 _07579_/S vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14139__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07836__A0 _15349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11632__A1 _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10435__A2 _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09240__B _15484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ _07486_/A vssd1 vssd1 vccd1 vccd1 _15521_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08137__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09225_ _15495_/Q vssd1 vssd1 vccd1 vccd1 _09225_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13978__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _09152_/A _09151_/B _09151_/A vssd1 vssd1 vccd1 vccd1 _09157_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__13697__B _13827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_884 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ _08107_/A vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__inv_2
XFILLER_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09087_ _15498_/Q _15482_/Q vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_110_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15771_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _12178_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08041_/B sky130_fd_sc_hd__xnor2_1
XFILLER_101_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14602__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _14934_/D sky130_fd_sc_hd__xor2_1
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09989_ _09990_/A _09990_/C _09990_/B vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__a21oi_1
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12122__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input139_A x_r_0[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _12426_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__nor2_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11961__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902_ _10902_/A _11117_/A _10902_/C vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__or3_1
X_11882_ _11882_/A _11963_/B vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__xnor2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14670_/Y sky130_fd_sc_hd__inv_2
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10833_ _15308_/Q _15143_/Q vssd1 vssd1 vccd1 vccd1 _10834_/C sky130_fd_sc_hd__and2b_1
XFILLER_83_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13621_ _15376_/Q _15360_/Q _13620_/B vssd1 vssd1 vccd1 vccd1 _13622_/B sky130_fd_sc_hd__a21o_1
XFILLER_198_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14049__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10764_ _15719_/Q _15785_/Q vssd1 vssd1 vccd1 vccd1 _10766_/A sky130_fd_sc_hd__or2b_1
X_13552_ _13552_/A _13552_/B vssd1 vssd1 vccd1 vccd1 _15600_/D sky130_fd_sc_hd__xnor2_1
XFILLER_197_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _14952_/Q _12510_/B vssd1 vssd1 vccd1 vccd1 _12614_/A sky130_fd_sc_hd__xnor2_2
XFILLER_13_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13483_ _13771_/B vssd1 vssd1 vccd1 vccd1 _13483_/Y sky130_fd_sc_hd__inv_2
X_10695_ _15280_/Q _15181_/Q vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0_1_clk clkbuf_1_0_1_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_199_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12434_ _12435_/A _12435_/B _12597_/A vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__o21ba_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15222_ _15498_/CLK _15222_/D _14270_/Y vssd1 vssd1 vccd1 vccd1 _15222_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12365_ _14940_/Q vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__inv_2
X_15153_ _15803_/CLK _15153_/D _14196_/Y vssd1 vssd1 vccd1 vccd1 _15153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_101_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15758_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11201__A _15028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14104_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14104_/Y sky130_fd_sc_hd__inv_2
X_11316_ _11317_/A _11317_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__xor2_1
XFILLER_10_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15084_ _15345_/CLK _15084_/D _14124_/Y vssd1 vssd1 vccd1 vccd1 _15084_/Q sky130_fd_sc_hd__dfrtp_1
X_12296_ _15739_/Q _12304_/B vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__and2_1
XANTENNA_output260_A _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output358_A _15682_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14035_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14035_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _11247_/A _11391_/A vssd1 vssd1 vccd1 vccd1 _11247_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14512__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ _15748_/Q _15026_/Q vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output525_A output525/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _10823_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _15798_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14937_ _15508_/CLK _14937_/D _13968_/Y vssd1 vssd1 vccd1 vccd1 _14937_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14868_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14868_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09118__B_N _15504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11590__B _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ _13819_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _15664_/D sky130_fd_sc_hd__xnor2_1
XFILLER_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14799_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14799_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09060__B _15364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_946 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09010_ _15371_/Q _15355_/Q vssd1 vssd1 vccd1 vccd1 _09010_/X sky130_fd_sc_hd__and2b_1
XFILLER_176_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09912_ _09983_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _14961_/D sky130_fd_sc_hd__xor2_1
XFILLER_160_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14422__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09843_ _15094_/Q vssd1 vssd1 vccd1 vccd1 _09843_/Y sky130_fd_sc_hd__inv_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _15429_/Q _15413_/Q _09772_/B _09773_/X vssd1 vssd1 vccd1 vccd1 _09775_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08725_ _08725_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _08725_/X sky130_fd_sc_hd__or2b_1
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08656_ _12644_/A _12644_/B vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__xor2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07607_ _07607_/A vssd1 vssd1 vccd1 vccd1 _15462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08587_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08711_/B sky130_fd_sc_hd__xor2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _15495_/Q input107/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07469_ _15529_/Q input93/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_69_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__A1 _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _09208_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _15298_/D sky130_fd_sc_hd__xor2_1
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _14901_/D sky130_fd_sc_hd__xor2_1
XFILLER_120_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_112_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ _15507_/Q _15491_/Q _09138_/X vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _12150_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12216_/B sky130_fd_sc_hd__xnor2_2
XFILLER_159_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11101_ _14936_/Q _15002_/Q vssd1 vssd1 vccd1 vccd1 _11101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11956__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _11997_/A _11997_/B _11994_/X vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__a21o_1
XFILLER_150_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_127_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14332__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input256_A x_r_7[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _14925_/Q _14991_/Q vssd1 vssd1 vccd1 vccd1 _11032_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08330__A _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13890__B _13890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15771_/CLK _15771_/D _14850_/Y vssd1 vssd1 vccd1 vccd1 _15771_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12981_/A _13547_/A _12982_/Y vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__o21ai_1
XFILLER_79_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11691__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14737_/A sky130_fd_sc_hd__buf_6
XFILLER_205_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11934_ _11867_/A _11867_/B _11868_/A vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__a21o_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09161__A _15566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14653_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11643_/A _11865_/B _11865_/C vssd1 vssd1 vccd1 vccd1 _11866_/D sky130_fd_sc_hd__and3b_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13604_ _15370_/Q _15354_/Q _13603_/X vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__a21oi_1
X_10816_ _10814_/A _10814_/B _10815_/X vssd1 vssd1 vccd1 vccd1 _10817_/B sky130_fd_sc_hd__a21o_1
X_11796_ _11796_/A _11777_/B vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__or2b_1
XFILLER_14_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14584_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14584_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _15760_/Q _13535_/B vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__nand2_1
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _10741_/A _10743_/B _10741_/B vssd1 vssd1 vccd1 vccd1 _10748_/B sky130_fd_sc_hd__a21boi_1
XFILLER_203_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14507__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13411__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10678_ _15276_/Q _15177_/Q _10674_/B vssd1 vssd1 vccd1 vccd1 _10679_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13466_ _13354_/A _13417_/A _13417_/B _13352_/A vssd1 vssd1 vccd1 vccd1 _13468_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output475_A output475/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ _15367_/CLK _15205_/D _14252_/Y vssd1 vssd1 vccd1 vccd1 _15205_/Q sky130_fd_sc_hd__dfrtp_1
X_12417_ _12416_/A _12455_/D _12455_/A vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__o21a_1
XFILLER_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13397_ _13443_/B _13397_/B vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__nor2_2
XFILLER_127_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _15400_/CLK _15136_/D _14178_/Y vssd1 vssd1 vccd1 vccd1 _15136_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12348_ _12332_/A _12331_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12348_/X sky130_fd_sc_hd__a21bo_1
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12279_ _12241_/B _12243_/B _12239_/Y vssd1 vssd1 vccd1 vccd1 _12280_/B sky130_fd_sc_hd__a21oi_2
X_15067_ _15346_/CLK _15067_/D _14106_/Y vssd1 vssd1 vccd1 vccd1 _15067_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14242__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07555__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14018_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14029_/A sky130_fd_sc_hd__buf_8
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08240__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater792_A _15601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08510_ _08504_/A _08504_/B _08509_/Y vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__a21oi_1
X_09490_ _15539_/Q vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08441_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08464_/A sky130_fd_sc_hd__xnor2_2
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_682 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _08396_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14417__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14152__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07465__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13991__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _15746_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09757_ _15067_/Q _15100_/Q vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__and2b_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _08713_/B vssd1 vssd1 vccd1 vccd1 _08709_/B sky130_fd_sc_hd__inv_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _15053_/Q vssd1 vssd1 vccd1 vccd1 _09688_/Y sky130_fd_sc_hd__inv_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ _08639_/A _08639_/B vssd1 vssd1 vccd1 vccd1 _08663_/B sky130_fd_sc_hd__and2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15133__D _15133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11506_/X _11501_/B _11576_/A _11576_/B _11507_/X vssd1 vssd1 vccd1 vccd1
+ _11651_/B sky130_fd_sc_hd__a221o_2
XFILLER_159_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _10519_/Y _10600_/B _10521_/B vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__o21ai_1
X_11581_ _15728_/Q _11581_/B vssd1 vssd1 vccd1 vccd1 _11581_/X sky130_fd_sc_hd__and2_1
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14972__D _14972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14327__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _13320_/A _13321_/A _13320_/C vssd1 vssd1 vccd1 vccd1 _13374_/A sky130_fd_sc_hd__or3_1
XFILLER_10_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10532_ _15259_/Q _15292_/Q vssd1 vssd1 vccd1 vccd1 _10532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ _10463_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _14896_/D sky130_fd_sc_hd__nor2_1
X_13251_ _13352_/A _15051_/Q _15052_/Q vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__and3_1
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ _12256_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__and2_1
X_13182_ _13255_/A _13182_/B vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__or2_1
X_10394_ _15106_/Q _15205_/Q vssd1 vssd1 vccd1 vccd1 _10395_/C sky130_fd_sc_hd__and2b_1
XANTENNA_input67_A x_i_4[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12133_ _12133_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__xor2_1
XFILLER_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07430__A1 _07430_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14062__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12064_ _12064_/A _12064_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__or2_1
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _11014_/A _11014_/B _10712_/B vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13109__C _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11625__S _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15754_/CLK _15754_/D _14832_/Y vssd1 vssd1 vccd1 vccd1 _15754_/Q sky130_fd_sc_hd__dfrtp_1
X_12966_ _12967_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__or2_1
XFILLER_166_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14705_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14705_/Y sky130_fd_sc_hd__inv_2
X_11917_ _11917_/A _11917_/B vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__xnor2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _15689_/CLK _15685_/D _14759_/Y vssd1 vssd1 vccd1 vccd1 _15685_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12897_/A _12923_/C vssd1 vssd1 vccd1 vccd1 _12940_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__15043__D _15043_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14636_/Y sky130_fd_sc_hd__inv_2
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11852_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10765__A _15785_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14567_/Y sky130_fd_sc_hd__inv_2
X_11779_ _11825_/B _11779_/B vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__xor2_4
XANTENNA__14237__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13518_ _13516_/Y _13588_/B _13515_/A _13514_/B _13517_/X vssd1 vssd1 vccd1 vccd1
+ _13527_/A sky130_fd_sc_hd__o221a_1
XFILLER_174_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14498_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater805_A _15584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13449_ _15770_/Q _13451_/A vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__xnor2_2
XFILLER_174_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15119_ _15119_/CLK _15119_/D _14161_/Y vssd1 vssd1 vccd1 vccd1 _15119_/Q sky130_fd_sc_hd__dfrtp_2
X_08990_ _15367_/Q vssd1 vssd1 vccd1 vccd1 _08990_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _10014_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _14938_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _15331_/Q _07872_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14700__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ _09611_/A _09611_/B _09806_/A vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__and3_1
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09542_ _15429_/Q _09542_/B _09772_/B vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__and3_1
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09473_ _09473_/A _09473_/B _09526_/A vssd1 vssd1 vccd1 vccd1 _09473_/X sky130_fd_sc_hd__and3_1
XFILLER_93_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08129__B _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15345_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08424_ _12654_/A _08396_/C _08423_/Y vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08355_ _15039_/Q vssd1 vssd1 vccd1 vccd1 _12810_/A sky130_fd_sc_hd__buf_6
XANTENNA__10675__A _15277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14147__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08286_ _08286_/A _08327_/A vssd1 vssd1 vccd1 vccd1 _08328_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08145__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13986__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07984__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07412__A1 _07412_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15128__D _15128_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14610__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ _09809_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _15166_/D sky130_fd_sc_hd__xnor2_1
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ _12820_/A _12820_/B vssd1 vssd1 vccd1 vccd1 _12826_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12130__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input121_A x_i_7[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input219_A x_r_5[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07479__A1 _07479_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ _12679_/A _12679_/B _12750_/Y vssd1 vssd1 vccd1 vccd1 _12800_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_81_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15791_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11702_ _11702_/A _11734_/C vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__xnor2_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15558_/CLK _15470_/D _14532_/Y vssd1 vssd1 vccd1 vccd1 _15470_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12755_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__xor2_1
XFILLER_163_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12784__B _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15798__D _15798_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14421_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14421_/Y sky130_fd_sc_hd__inv_2
X_11633_ _11633_/A _11633_/B vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__nor2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14057__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14352_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14352_/Y sky130_fd_sc_hd__inv_2
X_11564_ _11564_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__or2_1
XFILLER_210_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13303_ _15052_/Q _13303_/B vssd1 vssd1 vccd1 vccd1 _13350_/C sky130_fd_sc_hd__nor2_1
XFILLER_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07651__A1 _07651_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10598_/A sky130_fd_sc_hd__nand2_1
X_11495_ _11866_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11496_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14283_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10446_ _10445_/B _10445_/C _10445_/A vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__a21oi_1
X_13234_ _13234_/A _13333_/A vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _10375_/A _10484_/A _10376_/Y vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__o21ai_1
X_13165_ _13165_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__or2_1
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12041_/A _12041_/B _12040_/A vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__a21oi_1
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output340_A output340/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13096_ _13096_/A vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__inv_2
XFILLER_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15038__D _15038_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output438_A output438/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _12119_/A _12047_/B vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_914 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14520__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ _15808_/CLK _15806_/D _14886_/Y vssd1 vssd1 vccd1 vccd1 _15806_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_76 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13998_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14003_/A sky130_fd_sc_hd__buf_6
XFILLER_19_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15737_ _15790_/CLK _15737_/D _14814_/Y vssd1 vssd1 vccd1 vccd1 _15737_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12949_ _12949_/A _12870_/A vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__or2b_1
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater755_A repeater756/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 _15617_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15668_ _15670_/CLK _15668_/D _14741_/Y vssd1 vssd1 vccd1 vccd1 _15668_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_14619_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14619_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07890__A1 _07890_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater922_A repeater923/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _15705_/CLK _15599_/D _14669_/Y vssd1 vssd1 vccd1 vccd1 _15599_/Q sky130_fd_sc_hd__dfrtp_2
X_08140_ _11491_/A _08154_/B _08155_/B vssd1 vssd1 vccd1 vccd1 _08140_/X sky130_fd_sc_hd__or3_1
XFILLER_144_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08071_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08071_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07642__A1 _07642_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12215__A _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08973_ _08973_/A _08973_/B vssd1 vssd1 vccd1 vccd1 _15199_/D sky130_fd_sc_hd__xnor2_1
XFILLER_130_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07924_ _15561_/Q _15541_/Q vssd1 vssd1 vccd1 vccd1 _15284_/D sky130_fd_sc_hd__xor2_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14430__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07855_ _07855_/A vssd1 vssd1 vccd1 vccd1 _15340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13046__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _07786_/A vssd1 vssd1 vccd1 vccd1 _15374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09525_ _15536_/Q _15520_/Q _09524_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15690_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09456_ _15519_/Q _15535_/Q vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__or2b_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09870__A2 _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__nand2_2
XFILLER_61_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09387_ _09386_/A _09386_/C _09386_/B vssd1 vssd1 vccd1 vccd1 _09390_/C sky130_fd_sc_hd__a21o_1
XFILLER_196_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ _08329_/X _08292_/Y _08327_/X _08285_/Y _08337_/X vssd1 vssd1 vccd1 vccd1
+ _08338_/X sky130_fd_sc_hd__o221a_1
XFILLER_123_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12109__B _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08269_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__xor2_2
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14605__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ _10298_/Y _10300_/B vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__and2b_1
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ _11281_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11280_/X sky130_fd_sc_hd__xor2_4
XANTENNA__08603__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _15240_/Q vssd1 vssd1 vccd1 vccd1 _10231_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input169_A x_r_2[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10162_ _10160_/X _10168_/A vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput390 _15696_/Q vssd1 vssd1 vccd1 vccd1 y_i_7[4] sky130_fd_sc_hd__buf_2
XANTENNA__09138__A1 _15507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14970_ _15352_/CLK _14970_/D _14003_/Y vssd1 vssd1 vccd1 vccd1 _14970_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__nor2_2
XANTENNA__14340__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07653__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09153__B _15544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ _13728_/A _13732_/C _13837_/A vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _12803_/A _12803_/B vssd1 vssd1 vccd1 vccd1 _12805_/C sky130_fd_sc_hd__xnor2_1
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13783_ _13783_/A _13783_/B vssd1 vssd1 vccd1 vccd1 _13783_/X sky130_fd_sc_hd__or2_1
XFILLER_204_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10995_ _10994_/B _10994_/C _10994_/A vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_54_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15775_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15528_/CLK _15522_/D _14587_/Y vssd1 vssd1 vccd1 vccd1 _15522_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12996__A2 _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ _13022_/A _13022_/B _12733_/B vssd1 vssd1 vccd1 vccd1 _12777_/B sky130_fd_sc_hd__a21o_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07872__A1 _07872_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15453_ _15727_/CLK _15453_/D _14514_/Y vssd1 vssd1 vccd1 vccd1 _15453_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _12780_/A _12688_/A vssd1 vssd1 vccd1 vccd1 _12735_/B sky130_fd_sc_hd__nand2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14404_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14404_/Y sky130_fd_sc_hd__inv_2
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__or2_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _15803_/CLK _15384_/D _14442_/Y vssd1 vssd1 vccd1 vccd1 _15384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output290_A output290/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ _12596_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_560 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output388_A _15694_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__A1 _07624_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14335_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14335_/Y sky130_fd_sc_hd__inv_2
X_11547_ _11832_/A vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__inv_2
XFILLER_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14515__A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07828__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _14269_/A vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__inv_2
X_11478_ _11906_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08513__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_952 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13217_ _13217_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13217_/Y sky130_fd_sc_hd__nor2_1
X_10429_ _10428_/A _10428_/B _10078_/B vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__a21o_1
XFILLER_174_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14197_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14197_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ _13491_/S _14920_/Q vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__and2_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13079_ _13273_/A _13201_/A _13203_/A vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__and3b_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14250__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__B _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater872_A input256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07640_ _15445_/Q _07640_/A1 _07640_/S vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ _15479_/Q input43/X _07575_/S vssd1 vssd1 vccd1 vccd1 _07572_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15437_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_206_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ _09375_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _15127_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ _09239_/A _09239_/B _09240_/X vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__a21o_1
XFILLER_181_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09172_ _09170_/Y _09172_/B vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__nand2b_1
XFILLER_187_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ _08123_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__xor2_4
XFILLER_147_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14425__A _14439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ _12122_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08058_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07738__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08423__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput107 x_i_6[2] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_1
Xinput118 x_i_7[12] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07981__B _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14160__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _08882_/Y _08955_/B _08884_/B vssd1 vssd1 vccd1 vccd1 _08958_/B sky130_fd_sc_hd__o21ai_1
Xinput129 x_i_7[8] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07473__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07907_ _15461_/Q _15445_/Q vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__or2_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08887_ _08955_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _15209_/D sky130_fd_sc_hd__xor2_1
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater860 input42/X vssd1 vssd1 vccd1 vccd1 _07573_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater871 input3/X vssd1 vssd1 vccd1 vccd1 _07640_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ _15348_/Q input201/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07839_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater882 input244/X vssd1 vssd1 vccd1 vccd1 _07653_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater893 input230/X vssd1 vssd1 vccd1 vccd1 _07779_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07769_ _15382_/Q input154/X _07791_/S vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15433_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _15530_/Q _15514_/Q _09507_/X vssd1 vssd1 vccd1 vccd1 _09509_/B sky130_fd_sc_hd__a21oi_1
XFILLER_169_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10779_/A _10779_/B _11292_/A vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__a21o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07854__A1 input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09509_/A _09436_/B _09438_/X vssd1 vssd1 vccd1 vccd1 _09440_/B sky130_fd_sc_hd__a21o_1
XFILLER_200_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12450_ _14948_/Q vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__inv_2
XFILLER_8_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11401_ _10216_/A _11400_/B _10216_/B vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__14980__D _14980_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__A1 _07606_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12381_/A _12381_/B _12381_/C _12381_/D vssd1 vssd1 vccd1 vccd1 _12389_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14335__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14120_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11332_ _11333_/A _11333_/B vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__xor2_4
XFILLER_197_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14051_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11263_ _15713_/Q _11262_/Y _11261_/B vssd1 vssd1 vccd1 vccd1 _11265_/B sky130_fd_sc_hd__a21o_1
XFILLER_181_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__xnor2_1
XFILLER_180_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10214_ _15074_/Q _15239_/Q vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__or2_1
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11194_ _15027_/Q _15749_/Q vssd1 vssd1 vccd1 vccd1 _11195_/C sky130_fd_sc_hd__or2b_1
XFILLER_97_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10145_ _15145_/Q _15310_/Q vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__or2b_1
XFILLER_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14070__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14953_ _15784_/CLK _14953_/D _13985_/Y vssd1 vssd1 vccd1 vccd1 _14953_/Q sky130_fd_sc_hd__dfrtp_1
X_10076_ _15214_/Q _15115_/Q vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__and2b_1
XFILLER_47_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13904_ _15344_/Q _15328_/Q _13903_/B vssd1 vssd1 vccd1 vccd1 _13905_/B sky130_fd_sc_hd__a21o_1
XFILLER_208_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14884_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14884_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _14978_/Q vssd1 vssd1 vccd1 vccd1 _13836_/A sky130_fd_sc_hd__clkinv_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output303_A output303/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15399_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13414__A _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13766_ _14982_/Q _13858_/B vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__xnor2_2
X_10978_ _15271_/Q _10977_/Y _10976_/B vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15511_/CLK _15505_/D _14569_/Y vssd1 vssd1 vccd1 vccd1 _15505_/Q sky130_fd_sc_hd__dfrtp_4
X_12717_ _12717_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _12811_/A sky130_fd_sc_hd__xor2_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15051__D _15051_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ _14976_/Q _13827_/B vssd1 vssd1 vccd1 vccd1 _13826_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15436_ _15732_/CLK _15436_/D _14496_/Y vssd1 vssd1 vccd1 vccd1 _15436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__and2_1
XFILLER_54_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11869__A _12415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15367_ _15367_/CLK _15367_/D _14423_/Y vssd1 vssd1 vccd1 vccd1 _15367_/Q sky130_fd_sc_hd__dfrtp_2
X_12579_ _14940_/Q _12580_/B vssd1 vssd1 vccd1 vccd1 _12579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14245__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14318_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14318_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15298_ _15572_/CLK _15298_/D _14350_/Y vssd1 vssd1 vccd1 vccd1 _15298_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14249_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14249_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08810_/A _08818_/A vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__nand2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09790_ _15436_/Q _15420_/Q _09789_/X vssd1 vssd1 vccd1 vccd1 _09791_/B sky130_fd_sc_hd__a21oi_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__A0 _15376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__A _15495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08724_/X _08725_/X _08739_/X _08740_/X vssd1 vssd1 vccd1 vccd1 _08741_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08672_ _12688_/A _08672_/B _08672_/C vssd1 vssd1 vccd1 vccd1 _08672_/X sky130_fd_sc_hd__or3_1
XFILLER_113_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07623_ _07623_/A vssd1 vssd1 vccd1 vccd1 _15454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10948__A _10948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15749_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07554_ _07554_/A vssd1 vssd1 vccd1 vccd1 _15488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07485_ _15521_/Q input22/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07486_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _09224_/A _09224_/B vssd1 vssd1 vccd1 vccd1 _15236_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ _09153_/Y _09155_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__10683__A _15278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14155__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08106_ _08328_/A _08327_/A vssd1 vssd1 vccd1 vccd1 _08107_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09086_ _15498_/Q _15482_/Q vssd1 vssd1 vccd1 vccd1 _09086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13994__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08037_ _12122_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08041_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _15194_/Q _15227_/Q _09987_/B vssd1 vssd1 vccd1 vccd1 _09990_/C sky130_fd_sc_hd__a21o_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08939_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _15187_/D sky130_fd_sc_hd__xnor2_1
XFILLER_190_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09513__A1 _15532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _11950_/A _11950_/B vssd1 vssd1 vccd1 vccd1 _12022_/B sky130_fd_sc_hd__or2_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ _14894_/Q _14960_/Q vssd1 vssd1 vccd1 vccd1 _10902_/C sky130_fd_sc_hd__and2b_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater690 _14029_/A vssd1 vssd1 vccd1 vccd1 _14037_/A sky130_fd_sc_hd__buf_6
XFILLER_199_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11961__B _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14975__D _14975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _11957_/A _11881_/B vssd1 vssd1 vccd1 vccd1 _11963_/B sky130_fd_sc_hd__and2_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _13620_/A _13620_/B vssd1 vssd1 vccd1 vccd1 _15097_/D sky130_fd_sc_hd__nor2_1
X_10832_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__and2_1
XANTENNA_input201_A x_r_4[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__B _15515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13551_ _13551_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13552_/B sky130_fd_sc_hd__nor2_1
X_10763_ _11281_/A _10763_/B vssd1 vssd1 vccd1 vccd1 _10763_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_201_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12502_ _12502_/A _12502_/B vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__xor2_2
XFILLER_12_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13482_ _13477_/B _15771_/Q vssd1 vssd1 vccd1 vccd1 _13499_/B sky130_fd_sc_hd__and2b_1
XANTENNA_input97_A x_i_5[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ _15279_/Q _15180_/Q vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_699 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15221_ _15221_/CLK _15221_/D _14269_/Y vssd1 vssd1 vccd1 vccd1 _15221_/Q sky130_fd_sc_hd__dfrtp_1
X_12433_ _12431_/X _12433_/B vssd1 vssd1 vccd1 vccd1 _12597_/A sky130_fd_sc_hd__and2b_1
XFILLER_205_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14065__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _15170_/CLK _15152_/D _14195_/Y vssd1 vssd1 vccd1 vccd1 _15152_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_154_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12364_/A _12578_/A vssd1 vssd1 vccd1 vccd1 _15645_/D sky130_fd_sc_hd__xor2_1
XFILLER_165_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14103_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14103_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ _14925_/Q _11314_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _11317_/B sky130_fd_sc_hd__a21o_1
X_15083_ _15758_/CLK _15083_/D _14123_/Y vssd1 vssd1 vccd1 vccd1 _15083_/Q sky130_fd_sc_hd__dfrtp_4
X_12295_ _12493_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__xnor2_2
XFILLER_154_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14034_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _15758_/Q _15036_/Q vssd1 vssd1 vccd1 vccd1 _11391_/A sky130_fd_sc_hd__xnor2_2
XFILLER_180_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _15748_/Q _15026_/Q vssd1 vssd1 vccd1 vccd1 _11177_/Y sky130_fd_sc_hd__nor2_1
X_10128_ _10122_/A _10124_/B _10122_/B vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__a21boi_1
XANTENNA_output420_A output420/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15046__D _15046_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14936_ _15467_/CLK _14936_/D _13967_/Y vssd1 vssd1 vccd1 vccd1 _14936_/Q sky130_fd_sc_hd__dfrtp_2
X_10059_ _15210_/Q _15111_/Q _10055_/B vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__a21o_1
XFILLER_209_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14867_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14867_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater668_A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13818_ _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14798_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14798_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_550 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__A1 input178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _13748_/A _13748_/B _13748_/C vssd1 vssd1 vccd1 vccd1 _13849_/C sky130_fd_sc_hd__a21o_1
XANTENNA_repeater835_A input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ _15803_/CLK _15419_/D _14478_/Y vssd1 vssd1 vccd1 vccd1 _15419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11378__A1 _15753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12327__A0 _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14703__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _15191_/Q _09910_/Y _09906_/B vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09842_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _15750_/D sky130_fd_sc_hd__nor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13319__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _15430_/Q _15414_/Q vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__and2_1
XFILLER_6_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08622_/Y _08724_/B vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07506__A0 _15511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _13352_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07606_ _15462_/Q _07606_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08586_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__xor2_2
XFILLER_53_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13989__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ _07537_/A vssd1 vssd1 vccd1 vccd1 _15496_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12893__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07468_ _07468_/A vssd1 vssd1 vccd1 vccd1 _15530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09207_ _15575_/Q _15555_/Q vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07399_ _07399_/A vssd1 vssd1 vccd1 vccd1 _15568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09138_ _15507_/Q _15491_/Q _09133_/A vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09069_ _09222_/A _09069_/B vssd1 vssd1 vccd1 vccd1 _09219_/C sky130_fd_sc_hd__nand2_1
XFILLER_159_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14613__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11100_ _11100_/A _11350_/A vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__xor2_1
XFILLER_155_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12141_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11956__B _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11031_ _11309_/A _11031_/B vssd1 vssd1 vccd1 vccd1 _11031_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_78_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input151_A x_r_1[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input249_A x_r_7[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15770_ _15770_/CLK _15770_/D _14849_/Y vssd1 vssd1 vccd1 vccd1 _15770_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13294__A1 _13737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _15763_/Q _13549_/B vssd1 vssd1 vccd1 vccd1 _12982_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_894 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07661__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14721_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14721_/Y sky130_fd_sc_hd__inv_2
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A x_i_0[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11691__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__nand2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14652_/Y sky130_fd_sc_hd__inv_2
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _11710_/A _11861_/X _11866_/C _11712_/X _11863_/X vssd1 vssd1 vccd1 vccd1
+ _11867_/A sky130_fd_sc_hd__a221oi_2
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _15370_/Q _15354_/Q _13602_/B vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__o21a_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _15303_/Q _15138_/Q vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__and2b_1
XFILLER_60_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14583_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14583_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11795_ _11783_/A _11783_/B _11793_/X _11794_/X vssd1 vssd1 vccd1 vccd1 _11870_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_186_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _13534_/A vssd1 vssd1 vccd1 vccd1 _15596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10746_ _10744_/Y _10746_/B vssd1 vssd1 vccd1 vccd1 _11267_/A sky130_fd_sc_hd__and2b_1
XFILLER_199_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13465_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _10677_/A _11003_/A vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15204_ _15464_/CLK _15204_/D _14251_/Y vssd1 vssd1 vccd1 vccd1 _15204_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11212__A _11212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ _12416_/A _12455_/A _12455_/D vssd1 vssd1 vccd1 vccd1 _12418_/A sky130_fd_sc_hd__nor3_1
XFILLER_145_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output370_A output370/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _13396_/A _13396_/B _13396_/C vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__and3_1
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output468_A _11294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ _15400_/CLK _15135_/D _14177_/Y vssd1 vssd1 vccd1 vccd1 _15135_/Q sky130_fd_sc_hd__dfrtp_2
X_12347_ _15742_/Q _12522_/B vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__xor2_1
XFILLER_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14523__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07836__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15066_ _15346_/CLK _15066_/D _14105_/Y vssd1 vssd1 vccd1 vccd1 _15066_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12390__B_N _11728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12280_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08521__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10770__B _15785_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13139__A _13558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14017_/Y sky130_fd_sc_hd__inv_2
X_11229_ _11229_/A _11235_/A vssd1 vssd1 vccd1 vccd1 _11382_/A sky130_fd_sc_hd__nand2_2
XFILLER_136_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07571__S _07575_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater952_A input144/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ _15532_/CLK _14919_/D _13949_/Y vssd1 vssd1 vccd1 vccd1 _14919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08440_ _08459_/A _08458_/A vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__or2_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_694 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08404_/A sky130_fd_sc_hd__xor2_2
XFILLER_211_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08415__B _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__A1 _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14433__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11771__A1 _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A x_i_0[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _09824_/B _09824_/C _09824_/A vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__a21oi_1
XFILLER_154_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12888__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ _15066_/Q _15099_/Q vssd1 vssd1 vccd1 vccd1 _09760_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08707_ _08751_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _08707_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _15086_/Q _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nand2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__A1 _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08585_/X _08636_/Y _08637_/Y vssd1 vssd1 vccd1 vccd1 _08702_/A sky130_fd_sc_hd__a21bo_1
XFILLER_82_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08569_ _12662_/A vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__inv_2
XFILLER_202_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14608__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _14993_/D sky130_fd_sc_hd__xor2_1
X_11580_ _11580_/A _12529_/A vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__xor2_1
XFILLER_167_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_928 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ _10602_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__nand2_1
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input199_A x_r_4[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ _15051_/Q _13250_/B vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__nor2_1
XFILLER_182_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10462_ _10461_/B _10461_/C _10461_/A vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__a21oi_1
X_12201_ _12201_/A _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__nand3_1
XFILLER_164_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13181_ _13250_/B _13180_/C _13180_/A vssd1 vssd1 vccd1 vccd1 _13182_/B sky130_fd_sc_hd__o21a_1
XFILLER_164_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10393_ _10393_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _14942_/D sky130_fd_sc_hd__nor2_1
XFILLER_108_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14343__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _12204_/A _12131_/Y _12132_/S vssd1 vssd1 vccd1 vccd1 _12133_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09437__A _15532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12063_ _12063_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__or2_1
XFILLER_2_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _15019_/D sky130_fd_sc_hd__xor2_1
XFILLER_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _15754_/CLK _15753_/D _14831_/Y vssd1 vssd1 vccd1 vccd1 _15753_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _12965_/A _12965_/B vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__xor2_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11207__A _15030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ _12002_/B _11916_/B vssd1 vssd1 vccd1 vccd1 _11917_/B sky130_fd_sc_hd__xnor2_1
X_14704_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14704_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15684_ _15687_/CLK _15684_/D _14758_/Y vssd1 vssd1 vccd1 vccd1 _15684_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12896_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12923_/C sky130_fd_sc_hd__xor2_1
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14635_/Y sky130_fd_sc_hd__inv_2
X_11847_ _11908_/A _11907_/A vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__xor2_1
XFILLER_166_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13422__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14566_/Y sky130_fd_sc_hd__inv_2
X_11778_ _11797_/A _11797_/B vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__xnor2_2
XFILLER_186_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13517_ _13517_/A _13586_/A vssd1 vssd1 vccd1 vccd1 _13517_/X sky130_fd_sc_hd__or2b_1
XFILLER_53_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _15712_/Q _15778_/Q vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__or2_1
X_14497_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14497_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13448_ _13448_/A _13769_/B vssd1 vssd1 vccd1 vccd1 _13451_/A sky130_fd_sc_hd__xor2_2
XFILLER_70_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater700_A _07795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ _13431_/B _13379_/B vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14253__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15118_ _15367_/CLK _15118_/D _14160_/Y vssd1 vssd1 vccd1 vccd1 _15118_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_53_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08251__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _15086_/Q _15185_/Q vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__nor2_1
X_15049_ _15664_/CLK _15049_/D _14087_/Y vssd1 vssd1 vccd1 vccd1 _15049_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11505__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _07871_/A vssd1 vssd1 vccd1 vccd1 _15332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09610_ _09610_/A _09615_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__or2_1
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_68_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09541_ _15429_/Q _09542_/B _09772_/B vssd1 vssd1 vccd1 vccd1 _09545_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_111_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15812__A _15812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ _09472_/A _09480_/A vssd1 vssd1 vccd1 vccd1 _09526_/A sky130_fd_sc_hd__nand2_1
XFILLER_184_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10492__A1 _15251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08423_ _12810_/A _12654_/A vssd1 vssd1 vccd1 vccd1 _08423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14428__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_126_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08354_ _15726_/Q vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__inv_2
XFILLER_165_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08285_ _08288_/B _08285_/B vssd1 vssd1 vccd1 vccd1 _08285_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14163__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09257__A _09257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09808_ _09806_/A _09806_/B _09807_/X vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13226__B _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _09739_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__nand2_1
XFILLER_189_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ _12750_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _12750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input114_A x_i_6[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11701_ _11701_/A _11701_/B vssd1 vssd1 vccd1 vccd1 _11734_/C sky130_fd_sc_hd__xor2_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09720__A _15061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _08688_/A _08688_/B _12680_/Y vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14338__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14420_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14439_/A sky130_fd_sc_hd__buf_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _12244_/A _11631_/B _11631_/C vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__a21oi_1
XFILLER_187_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14351_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14351_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ _11563_/A vssd1 vssd1 vccd1 vccd1 _11563_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _15052_/Q _13303_/B vssd1 vssd1 vccd1 vccd1 _13356_/A sky130_fd_sc_hd__and2_1
XFILLER_155_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _15256_/Q _15289_/Q vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14282_/Y sky130_fd_sc_hd__inv_2
X_11494_ _11493_/A _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11697__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ _13233_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13333_/A sky130_fd_sc_hd__and2_1
XFILLER_183_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _10445_/A _10445_/B _10445_/C vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__and3_1
XFILLER_100_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14073__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07386__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13164_ _13222_/A _13222_/B vssd1 vssd1 vccd1 vccd1 _13219_/A sky130_fd_sc_hd__xnor2_1
X_10376_ _15134_/Q _15167_/Q vssd1 vssd1 vccd1 vccd1 _10376_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12115_ _12160_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13095_ _13097_/A _13097_/B _13097_/C vssd1 vssd1 vccd1 vccd1 _13096_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__14801__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12046_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12047_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output333_A _11348_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15805_ _15808_/CLK _15805_/D _14885_/Y vssd1 vssd1 vccd1 vccd1 _15805_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13997_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13997_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15736_ _15790_/CLK _15736_/D _14813_/Y vssd1 vssd1 vccd1 vccd1 _15736_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__A1 _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ _12985_/C _12985_/B _13020_/B vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__a21o_1
XFILLER_46_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater650_A _07971_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ _15680_/CLK _15667_/D _14740_/Y vssd1 vssd1 vccd1 vccd1 _15667_/Q sky130_fd_sc_hd__dfrtp_1
X_12879_ _13021_/A _13021_/B _13022_/B _13022_/A vssd1 vssd1 vccd1 vccd1 _12909_/B
+ sky130_fd_sc_hd__or4bb_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater748_A _15654_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14248__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14618_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14618_/Y sky130_fd_sc_hd__inv_2
X_15598_ _15707_/CLK _15598_/D _14668_/Y vssd1 vssd1 vccd1 vccd1 _15598_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08246__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14549_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14549_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater915_A input198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ _08070_/A _08070_/B vssd1 vssd1 vccd1 vccd1 _08086_/A sky130_fd_sc_hd__xnor2_2
XFILLER_146_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08972_ _08970_/A _08970_/B _08971_/X vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14711__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07923_ _07923_/A vssd1 vssd1 vccd1 vccd1 _15152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13327__A _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07854_ _15340_/Q input208/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12231__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07785_ _15374_/Q _07785_/A1 _07803_/S vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__mux2_1
XFILLER_209_280 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _15262_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10465__A1 _15127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09455_ _15534_/Q _15518_/Q vssd1 vssd1 vccd1 vccd1 _09459_/B sky130_fd_sc_hd__or2b_1
XFILLER_197_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10686__A _15278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14158__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _08392_/Y _08405_/A _08403_/X _08441_/B _08441_/A vssd1 vssd1 vccd1 vccd1
+ _08443_/B sky130_fd_sc_hd__a32o_1
XFILLER_197_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09386_ _09386_/A _09386_/B _09386_/C vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__and3_1
XFILLER_61_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08337_ _11678_/A _11545_/A _08329_/X _08292_/Y _08336_/X vssd1 vssd1 vccd1 vccd1
+ _08337_/X sky130_fd_sc_hd__a221o_1
XFILLER_196_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13997__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09428__A_N _15529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08268_ _08321_/A _08264_/Y _08273_/B _08273_/A vssd1 vssd1 vccd1 vccd1 _08269_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_193_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__or2b_1
XFILLER_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10230_ _10230_/A _10230_/B vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__nand2_2
XFILLER_133_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10161_ _10160_/A _10160_/B _10848_/A vssd1 vssd1 vccd1 vccd1 _10168_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput380 output380/A vssd1 vssd1 vccd1 vccd1 y_i_7[10] sky130_fd_sc_hd__buf_2
XFILLER_86_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput391 output391/A vssd1 vssd1 vccd1 vccd1 y_i_7[5] sky130_fd_sc_hd__buf_2
XFILLER_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09138__A2 _15491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14978__D _14978_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ _15117_/Q _15216_/Q vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__and2b_1
XFILLER_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input231_A x_r_6[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13920_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09434__B _15514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13851_ _13752_/A _13752_/B _13838_/C _13842_/A _13838_/B vssd1 vssd1 vccd1 vccd1
+ _13851_/X sky130_fd_sc_hd__o2111a_1
XFILLER_142_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12802_ _12802_/A _12872_/A vssd1 vssd1 vccd1 vccd1 _12803_/B sky130_fd_sc_hd__xnor2_1
X_13782_ _13792_/B _13782_/B vssd1 vssd1 vccd1 vccd1 _13785_/A sky130_fd_sc_hd__xnor2_1
X_10994_ _10994_/A _10994_/B _10994_/C vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__or3_1
XFILLER_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _13022_/A _12733_/B _13022_/B vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__nand3_1
X_15521_ _15532_/CLK _15521_/D _14586_/Y vssd1 vssd1 vccd1 vccd1 _15521_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14068__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15452_ _15558_/CLK _15452_/D _14513_/Y vssd1 vssd1 vccd1 vccd1 _15452_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_203_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12664_ _12780_/A _08675_/B _08677_/Y _12663_/Y vssd1 vssd1 vccd1 vccd1 _12683_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14403_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14403_/Y sky130_fd_sc_hd__inv_2
X_11615_ _11615_/A _11615_/B vssd1 vssd1 vccd1 vccd1 _12378_/B sky130_fd_sc_hd__xnor2_4
XFILLER_169_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ _15383_/CLK _15383_/D _14439_/Y vssd1 vssd1 vccd1 vccd1 _15383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12595_ _12420_/A _12425_/B _12593_/B _12593_/A vssd1 vssd1 vccd1 vccd1 _12596_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14334_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14334_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11546_ _11928_/A _11832_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11620_/B sky130_fd_sc_hd__and3_1
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output283_A _15658_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14265_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14265_/Y sky130_fd_sc_hd__inv_2
X_11477_ _11559_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09609__B _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A _15754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13216_ _13247_/B _13216_/B vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__and2_1
XFILLER_171_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _14951_/D sky130_fd_sc_hd__xor2_2
XANTENNA_output450_A output450/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14196_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07388__A1 _07388_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__B _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13147_/A _13147_/B vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__nand2_1
X_10359_ _10359_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__nor2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14531__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07844__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13265_/B _13078_/B vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__nor2_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater698_A _07795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12029_ _12029_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__or2b_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13881__A1 _15336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater865_A repeater866/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ _07570_/A vssd1 vssd1 vccd1 vccd1 _15480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15719_ _15719_/CLK _15719_/D _14795_/Y vssd1 vssd1 vccd1 vccd1 _15719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12987__A3 _12976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09240_ _15500_/Q _15484_/Q vssd1 vssd1 vccd1 vccd1 _09240_/X sky130_fd_sc_hd__and2b_1
XFILLER_146_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09171_ _15568_/Q _15548_/Q vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14706__A _14709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _08272_/A _08119_/Y _08271_/B _08271_/A vssd1 vssd1 vccd1 vccd1 _08123_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08704__A _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ _12055_/A _08077_/B vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__nand2_1
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08423__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 x_i_6[3] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_2
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08955_ _08955_/A _08955_/B vssd1 vssd1 vccd1 vccd1 _15193_/D sky130_fd_sc_hd__xor2_1
Xinput119 x_i_7[13] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12124__A1 _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07906_ _15461_/Q _15445_/Q vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__nand2_1
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08886_ _08952_/A _08881_/B _08885_/X vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater850 repeater851/X vssd1 vssd1 vccd1 vccd1 _07441_/A1 sky130_fd_sc_hd__buf_4
XFILLER_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater861 input41/X vssd1 vssd1 vccd1 vccd1 _07545_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07837_ _07837_/A vssd1 vssd1 vccd1 vccd1 _15349_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A1 _07551_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater872 input256/X vssd1 vssd1 vccd1 vccd1 _07659_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13491__S _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater883 input242/X vssd1 vssd1 vccd1 vccd1 _07785_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater894 input228/X vssd1 vssd1 vccd1 vccd1 _07783_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07768_ _07768_/A vssd1 vssd1 vccd1 vccd1 _15383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09507_ _15530_/Q _15514_/Q _09506_/B vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07699_ _07699_/A vssd1 vssd1 vccd1 vccd1 _07750_/S sky130_fd_sc_hd__buf_12
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _15531_/Q _15515_/Q vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__and2b_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _15403_/Q _15387_/Q vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__and2b_1
XFILLER_166_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14616__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11400_ _11400_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _15731_/D sky130_fd_sc_hd__xnor2_2
X_12380_ _12381_/B _12381_/C _12381_/D _12381_/A vssd1 vssd1 vccd1 vccd1 _12391_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08614__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _14929_/Q _11330_/Y _11329_/B vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__a21o_1
XANTENNA_input181_A x_r_3[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08333__B _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14050_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14050_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11262_ _15779_/Q vssd1 vssd1 vccd1 vccd1 _11262_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _13201_/A _12714_/B _13000_/Y vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__a21oi_1
X_10213_ _10213_/A _10213_/B vssd1 vssd1 vccd1 vccd1 _15762_/D sky130_fd_sc_hd__nor2_1
XFILLER_134_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14351__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _11191_/Y _11193_/B vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__and2b_2
XANTENNA_input42_A x_i_2[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10834_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _15801_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _15784_/CLK _14952_/D _13984_/Y vssd1 vssd1 vccd1 vccd1 _14952_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ _15213_/Q _15114_/Q vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13903_ _13903_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _15064_/D sky130_fd_sc_hd__nor2_1
X_14883_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14883_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ _13838_/C _13834_/B vssd1 vssd1 vccd1 vccd1 _15668_/D sky130_fd_sc_hd__nor2_2
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11221__B_N _15754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _13772_/B _13765_/B vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__or2_1
X_10977_ _15172_/Q vssd1 vssd1 vccd1 vccd1 _10977_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15504_ _15511_/CLK _15504_/D _14568_/Y vssd1 vssd1 vccd1 vccd1 _15504_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_204_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _12827_/A _12827_/B vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__xor2_1
X_13696_ _13696_/A _13696_/B vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__xnor2_1
XFILLER_189_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ _15435_/CLK _15435_/D _14495_/Y vssd1 vssd1 vccd1 vccd1 _15435_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_175_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12647_ _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__nor2_1
XFILLER_203_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14526__A _14526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13430__A _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15366_ _15460_/CLK _15366_/D _14422_/Y vssd1 vssd1 vccd1 vccd1 _15366_/Q sky130_fd_sc_hd__dfrtp_1
X_12578_ _12578_/A _12578_/B vssd1 vssd1 vccd1 vccd1 _15678_/D sky130_fd_sc_hd__xor2_1
XFILLER_156_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _11585_/B _11529_/B vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__xnor2_1
XFILLER_141_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14317_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14317_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater613_A _10889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15297_ _15572_/CLK _15297_/D _14349_/Y vssd1 vssd1 vccd1 vccd1 _15297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14248_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14248_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14179_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14198_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_113_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14261__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater982_A input112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07781__A1 input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08621_/A _08621_/B _08624_/A vssd1 vssd1 vccd1 vccd1 _08740_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08671_ _08671_/A _08671_/B vssd1 vssd1 vccd1 vccd1 _13634_/A sky130_fd_sc_hd__xnor2_4
X_07622_ _15454_/Q input18/X _07644_/S vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07553_ _15488_/Q input37/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07554_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15242__D _15242_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07484_ _07484_/A vssd1 vssd1 vccd1 vccd1 _15522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _09222_/A _09222_/C _09222_/B vssd1 vssd1 vccd1 vccd1 _09224_/B sky130_fd_sc_hd__a21oi_2
XFILLER_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1097 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14436__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09154_ _15564_/Q _15544_/Q vssd1 vssd1 vccd1 vccd1 _09155_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08434__A _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08105_ _08105_/A _08105_/B _08329_/A vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__or3_1
X_09085_ _09230_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _15222_/D sky130_fd_sc_hd__xnor2_1
XFILLER_120_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08036_ _08036_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08054_/B sky130_fd_sc_hd__xnor2_1
XFILLER_163_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 x_i_5[1] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14171__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09987_ _09987_/A _09987_/B vssd1 vssd1 vccd1 vccd1 _14930_/D sky130_fd_sc_hd__xnor2_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__B _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08938_ _15461_/Q _15445_/Q _08936_/B _08937_/X vssd1 vssd1 vccd1 vccd1 _08939_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _15465_/Q _15449_/Q vssd1 vssd1 vccd1 vccd1 _08869_/X sky130_fd_sc_hd__and2b_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__A1 _07524_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__nand2_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater680 _14515_/A vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__buf_4
XFILLER_17_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ _12238_/A _12231_/A vssd1 vssd1 vccd1 vccd1 _11881_/B sky130_fd_sc_hd__or2_1
Xrepeater691 _14003_/A vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__buf_8
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _14912_/D sky130_fd_sc_hd__xor2_4
XFILLER_198_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _13549_/A _13549_/B _13546_/B _13546_/A vssd1 vssd1 vccd1 vccd1 _13551_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ _10754_/Y _10758_/B _10756_/B vssd1 vssd1 vccd1 vccd1 _10763_/B sky130_fd_sc_hd__o21ai_2
XFILLER_73_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _12500_/Y _12493_/B _12292_/B vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__a21o_1
XFILLER_186_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ _13499_/A _13481_/B vssd1 vssd1 vccd1 vccd1 _15639_/D sky130_fd_sc_hd__nor2_1
XFILLER_197_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ _10693_/A vssd1 vssd1 vccd1 vccd1 _15048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14346__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ _15220_/CLK _15220_/D _14268_/Y vssd1 vssd1 vccd1 vccd1 _15220_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13250__A _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _14946_/Q _12440_/C _12438_/B vssd1 vssd1 vccd1 vccd1 _12433_/B sky130_fd_sc_hd__or3_1
XANTENNA__07659__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15151_ _15394_/CLK _15151_/D _14194_/Y vssd1 vssd1 vccd1 vccd1 _15151_/Q sky130_fd_sc_hd__dfrtp_1
X_12363_ _14940_/Q _12580_/B vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__xnor2_2
XFILLER_181_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14102_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14102_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ _14991_/Q vssd1 vssd1 vccd1 vccd1 _11314_/Y sky130_fd_sc_hd__inv_2
X_15082_ _15758_/CLK _15082_/D _14122_/Y vssd1 vssd1 vccd1 vccd1 _15082_/Q sky130_fd_sc_hd__dfrtp_1
X_12294_ _12261_/X _12265_/B _12263_/B vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__o21ai_2
XFILLER_181_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14033_/Y sky130_fd_sc_hd__inv_2
X_11245_ _11243_/A _11388_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11247_/A sky130_fd_sc_hd__o21a_1
XFILLER_122_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14081__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07394__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11176_ _11361_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07763__A1 _07763_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10127_ _10125_/Y _10127_/B vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14935_ _15508_/CLK _14935_/D _13966_/Y vssd1 vssd1 vccd1 vccd1 _14935_/Q sky130_fd_sc_hd__dfrtp_2
X_10058_ _10058_/A _10421_/A vssd1 vssd1 vccd1 vccd1 _10417_/A sky130_fd_sc_hd__nand2_2
XFILLER_209_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output413_A output413/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14866_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08519__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13817_ _13816_/A _13816_/B _13812_/B _13812_/A _13813_/X vssd1 vssd1 vccd1 vccd1
+ _13818_/B sky130_fd_sc_hd__o221a_1
XFILLER_17_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater563_A _11134_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14797_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14797_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_904 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13748_ _13748_/A _13748_/B _13748_/C vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__nand3_1
XFILLER_91_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater730_A _15678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater828_A input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ _12985_/B _12910_/C _12910_/A vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__a21bo_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14256__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07569__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15418_ _15434_/CLK _15418_/D _14477_/Y vssd1 vssd1 vccd1 vccd1 _15418_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11378__A2 _15031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15349_ _15354_/CLK _15349_/D _14404_/Y vssd1 vssd1 vccd1 vccd1 _15349_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ _15224_/Q vssd1 vssd1 vccd1 vccd1 _09910_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _09840_/B _09840_/C _09840_/A vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15237__D _15237_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15815__A _15815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _09772_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _15153_/D sky130_fd_sc_hd__xnor2_1
XFILLER_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08723_ _12921_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _08723_/X sky130_fd_sc_hd__or2_1
XFILLER_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07506__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__xnor2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07605_ _07605_/A vssd1 vssd1 vccd1 vccd1 _15463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08751_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _08585_/X sky130_fd_sc_hd__or2_1
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07536_ _15496_/Q input108/X _07536_/S vssd1 vssd1 vccd1 vccd1 _07537_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12893__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07987__B _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ _15530_/Q _07467_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14166__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__A _15279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _09204_/A _09674_/A _09205_/Y vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07479__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08164__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07398_ _15568_/Q _07398_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07399_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09137_ _09137_/A vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_194_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ _15478_/Q _15494_/Q vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__or2b_1
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08019_ _11898_/A _11797_/A vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__xor2_2
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12414__A _14945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11030_ _11026_/A _11023_/Y _11025_/B vssd1 vssd1 vccd1 vccd1 _11031_/B sky130_fd_sc_hd__o21ai_2
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input144_A x_r_0[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _12981_/A _13547_/A vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__xor2_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14720_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14720_/Y sky130_fd_sc_hd__inv_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11932_ _11932_/A vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__inv_2
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11863_ _11753_/B _11863_/B vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__and2b_1
X_14651_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10814_/A _10814_/B vssd1 vssd1 vccd1 vccd1 _14907_/D sky130_fd_sc_hd__xor2_1
X_13602_ _13602_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _15091_/D sky130_fd_sc_hd__xnor2_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _12403_/B _12403_/A vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__or2b_1
X_14582_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14582_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10745_ _15715_/Q _15781_/Q vssd1 vssd1 vccd1 vccd1 _10746_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13533_ _13536_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__and2_1
XFILLER_198_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14076__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07681__A0 _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ _13464_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__xnor2_4
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08074__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _15178_/Q _15277_/Q vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__or2b_1
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_83 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12415_ _11938_/B _12415_/B vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__and2b_1
XFILLER_12_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15203_ _15464_/CLK _15203_/D _14250_/Y vssd1 vssd1 vccd1 vccd1 _15203_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _13396_/A _13396_/B _13396_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14804__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _12346_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__xnor2_2
XFILLER_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15134_ _15428_/CLK _15134_/D _14176_/Y vssd1 vssd1 vccd1 vccd1 _15134_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output363_A output363/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _15758_/CLK _15065_/D _14104_/Y vssd1 vssd1 vccd1 vccd1 _15065_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_494 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12277_ _12277_/A _12277_/B vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__or2_1
XFILLER_4_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14016_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14016_/Y sky130_fd_sc_hd__inv_2
X_11228_ _15033_/Q _15755_/Q vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__or2b_1
XANTENNA_output530_A output530/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07736__A1 input218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ _15022_/Q vssd1 vssd1 vccd1 vccd1 _11159_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07852__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater680_A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater778_A repeater779/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__A2 _13563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14918_ _15532_/CLK _14918_/D _13948_/Y vssd1 vssd1 vccd1 vccd1 _14918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14849_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12994__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater945_A input153/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _13273_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13602__B _13602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14714__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09824_ _09824_/A _09824_/B _09824_/C vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__and3_1
XFILLER_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12888__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09755_ _09755_/A vssd1 vssd1 vccd1 vccd1 _15722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08706_ _08706_/A vssd1 vssd1 vccd1 vccd1 _15594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _09686_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _15710_/D sky130_fd_sc_hd__xnor2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08637_ _08751_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _08637_/Y sky130_fd_sc_hd__nand2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13028__A2 _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07998__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _13046_/A vssd1 vssd1 vccd1 vccd1 _08570_/A sky130_fd_sc_hd__inv_2
XFILLER_39_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07519_ _07519_/A vssd1 vssd1 vccd1 vccd1 _15505_/D sky130_fd_sc_hd__clkbuf_1
X_08499_ _12803_/A _12688_/A _08499_/C vssd1 vssd1 vccd1 vccd1 _08508_/B sky130_fd_sc_hd__and3_1
XFILLER_211_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ _10602_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _15027_/D sky130_fd_sc_hd__xor2_1
XFILLER_156_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _10461_/A _10461_/B _10461_/C vssd1 vssd1 vccd1 vccd1 _10463_/A sky130_fd_sc_hd__and3_1
XFILLER_6_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13803__B_N _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14624__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12201_/A _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__a21o_1
XFILLER_182_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13180_ _13180_/A _13250_/B _13180_/C vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__nor3_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10392_ _10391_/B _10391_/C _10391_/A vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12131_ _12204_/A _12144_/A vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12144__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _12062_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__or2b_1
XFILLER_150_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07718__A1 input212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ _11012_/A _11012_/B _10705_/B vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15605__D _15605_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15752_/CLK _15752_/D _14830_/Y vssd1 vssd1 vccd1 vccd1 _15752_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _13046_/A _12858_/B _12863_/B _12963_/X vssd1 vssd1 vccd1 vccd1 _12965_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08069__A _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14703_/Y sky130_fd_sc_hd__inv_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11915_ _11991_/A _11697_/C _12088_/A vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15687_/CLK _15683_/D _14757_/Y vssd1 vssd1 vccd1 vccd1 _15683_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12937_/A _12937_/B vssd1 vssd1 vccd1 vccd1 _12896_/B sky130_fd_sc_hd__xnor2_1
XFILLER_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14634_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14634_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11846_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11907_/A sky130_fd_sc_hd__xnor2_1
XFILLER_127_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11777_ _11796_/A _11777_/B vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__xnor2_1
XFILLER_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14565_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14565_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10728_ _10728_/A _11251_/B vssd1 vssd1 vccd1 vccd1 _10728_/Y sky130_fd_sc_hd__xnor2_4
X_13516_ _15773_/Q vssd1 vssd1 vccd1 vccd1 _13516_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output480_A _11280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14496_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14496_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _10982_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _15042_/D sky130_fd_sc_hd__xnor2_4
X_13447_ _13770_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13769_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__14534__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09628__A _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__A1 _15750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _13433_/A _13378_/B vssd1 vssd1 vccd1 vccd1 _13379_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12950__A1 _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15117_ _15346_/CLK _15117_/D _14158_/Y vssd1 vssd1 vccd1 vccd1 _15117_/Q sky130_fd_sc_hd__dfrtp_1
X_12329_ _12329_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12330_/S sky130_fd_sc_hd__or2b_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08251__B _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ _15664_/CLK _15048_/D _14086_/Y vssd1 vssd1 vccd1 vccd1 _15048_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater895_A input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07870_ _15332_/Q _07870_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_478 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _09545_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__or2_1
XFILLER_3_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09471_ _15537_/Q _15521_/Q vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__or2b_1
XANTENNA__09882__A1 _15187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14709__A _14709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08422_ _12921_/A _12810_/A _08422_/C vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__and3_1
XFILLER_97_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ _08353_/A vssd1 vssd1 vccd1 vccd1 _15643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12229__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15250__D _15250_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ _11832_/A _08292_/B _08288_/A _08252_/D vssd1 vssd1 vccd1 vccd1 _08285_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14444__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07757__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08373__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07492__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09807_ _15442_/Q _15426_/Q vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__and2_1
XFILLER_8_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07999_ _15799_/Q vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__buf_6
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09738_ _09739_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _15720_/D sky130_fd_sc_hd__xor2_1
XANTENNA__13226__C _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09669_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _15312_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14619__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11746_/B _11700_/B vssd1 vssd1 vccd1 vccd1 _11701_/B sky130_fd_sc_hd__xor2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _12680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_203_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A x_i_6[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _12244_/A _11631_/B _11631_/C vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__and3_1
XFILLER_30_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07636__A0 _15447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11562_ _11562_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__xnor2_1
X_14350_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14350_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ _15256_/Q _15289_/Q vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__or2_1
X_13301_ _13301_/A _13301_/B vssd1 vssd1 vccd1 vccd1 _13303_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__inv_2
X_11493_ _11493_/A _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11866_/A sky130_fd_sc_hd__nand3_2
XFILLER_109_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14354__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07667__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ _13233_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13234_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11697__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10444_ _15155_/Q _15122_/Q vssd1 vssd1 vccd1 vccd1 _10445_/C sky130_fd_sc_hd__or2b_1
XANTENNA_input72_A x_i_4[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13163_ _13113_/A _13113_/B _13162_/X vssd1 vssd1 vccd1 vccd1 _13222_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10375_ _10375_/A _10484_/A vssd1 vssd1 vccd1 vccd1 _15790_/D sky130_fd_sc_hd__xor2_1
XFILLER_152_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12114_ _12167_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__and2_1
XFILLER_112_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ _13203_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _13097_/C sky130_fd_sc_hd__xnor2_1
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12045_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12119_/A sky130_fd_sc_hd__and2_1
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _15808_/CLK _15804_/D _14884_/Y vssd1 vssd1 vccd1 vccd1 _15804_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13996_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15735_ _15790_/CLK _15735_/D _14812_/Y vssd1 vssd1 vccd1 vccd1 _15735_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12947_ _12985_/C _12985_/B _13020_/B vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__nand3_1
XFILLER_18_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14529__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15666_ _15666_/CLK _15666_/D _14739_/Y vssd1 vssd1 vccd1 vccd1 _15666_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12973_/B _12878_/B vssd1 vssd1 vccd1 vccd1 _12910_/A sky130_fd_sc_hd__or2_2
XFILLER_60_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10776__B _15787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14617_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14617_/Y sky130_fd_sc_hd__inv_2
X_11829_ _11829_/A _11829_/B _11829_/C vssd1 vssd1 vccd1 vccd1 _11831_/A sky130_fd_sc_hd__nand3_1
XANTENNA_repeater643_A _11149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15597_ _15707_/CLK _15597_/D _14667_/Y vssd1 vssd1 vccd1 vccd1 _15597_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14548_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14548_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater810_A _15577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14479_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14479_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14264__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07577__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__A _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08971_ _15474_/Q _15458_/Q vssd1 vssd1 vccd1 vccd1 _08971_/X sky130_fd_sc_hd__and2_1
XFILLER_29_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07922_ _09772_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07923_/A sky130_fd_sc_hd__and2_1
XFILLER_190_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07853_ _07853_/A vssd1 vssd1 vccd1 vccd1 _15341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07784_ _07784_/A vssd1 vssd1 vccd1 vccd1 _15375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _09522_/B _09522_/C _09522_/A vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__o21a_1
XFILLER_209_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14439__A _14439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09454_ _09516_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08405_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08441_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13062__B _13062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _09385_/A vssd1 vssd1 vccd1 vccd1 _15145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07618__A0 _15456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _11678_/A _11545_/A _11480_/A _11658_/A _08335_/X vssd1 vssd1 vccd1 vccd1
+ _08336_/X sky130_fd_sc_hd__o221a_1
XFILLER_162_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08267_ _08267_/A vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__inv_2
XFILLER_20_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14174__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08198_ _11617_/A _11467_/A vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__nand2_1
XFILLER_180_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ _10160_/A _10160_/B _10848_/A vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__and3_1
XFILLER_161_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput370 output370/A vssd1 vssd1 vccd1 vccd1 y_i_6[1] sky130_fd_sc_hd__buf_2
XFILLER_160_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput381 output381/A vssd1 vssd1 vccd1 vccd1 y_i_7[11] sky130_fd_sc_hd__buf_2
XFILLER_156_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput392 _15698_/Q vssd1 vssd1 vccd1 vccd1 y_i_7[6] sky130_fd_sc_hd__buf_2
XFILLER_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ _15216_/Q _15117_/Q vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__and2b_1
XFILLER_48_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input224_A x_r_5[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ _13752_/A _13752_/B _13847_/A vssd1 vssd1 vccd1 vccd1 _13850_/X sky130_fd_sc_hd__o21ba_1
XFILLER_142_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _12799_/Y _12753_/B _12800_/Y vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__o21a_1
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10993_ _15176_/Q _15275_/Q vssd1 vssd1 vccd1 vccd1 _10994_/C sky130_fd_sc_hd__and2b_1
X_13781_ _13781_/A _13781_/B vssd1 vssd1 vccd1 vccd1 _13792_/B sky130_fd_sc_hd__and2_1
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14349__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13253__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _15563_/CLK _15520_/D _14585_/Y vssd1 vssd1 vccd1 vccd1 _15520_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _08671_/A _08671_/B _12657_/B _12658_/X vssd1 vssd1 vccd1 vccd1 _13022_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_203_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_615 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_52_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15553_/CLK _15451_/D _14512_/Y vssd1 vssd1 vccd1 vccd1 _15451_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12663_/Y sky130_fd_sc_hd__nand2_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14402_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14402_/Y sky130_fd_sc_hd__inv_2
X_11614_ _11828_/A _11827_/C _11828_/B _11538_/A vssd1 vssd1 vccd1 vccd1 _11615_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_187_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15382_ _15666_/CLK _15382_/D _14438_/Y vssd1 vssd1 vccd1 vccd1 _15382_/Q sky130_fd_sc_hd__dfrtp_1
X_12594_ _12594_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _15683_/D sky130_fd_sc_hd__xor2_1
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14333_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__inv_2
X_11545_ _11545_/A _11687_/A _11617_/A vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__and3_1
XFILLER_11_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_67_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14084__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15493_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11476_ _12247_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__xnor2_1
X_14264_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14264_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_110_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output276_A output276/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13215_ _15767_/Q vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__inv_2
X_10427_ _10426_/A _10426_/B _10070_/B vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__a21o_1
X_14195_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14195_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14812__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__C _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10358_ _15165_/Q _15132_/Q vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__and2b_1
X_13146_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13147_/B sky130_fd_sc_hd__inv_2
XFILLER_174_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output443_A output443/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13077_ _13352_/A _13366_/A _13076_/C vssd1 vssd1 vccd1 vccd1 _13078_/B sky130_fd_sc_hd__a21oi_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12332__A _12332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _10287_/A _11427_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10291_/A sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_125_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A1 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _12126_/A _12126_/B vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__nand2_2
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater593_A _10763_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07860__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater760_A _15642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13979_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14259__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15718_ _15719_/CLK _15718_/D _14794_/Y vssd1 vssd1 vccd1 vccd1 _15718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15649_ _15649_/CLK _15649_/D _14721_/Y vssd1 vssd1 vccd1 vccd1 _15649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _15568_/Q _15548_/Q vssd1 vssd1 vccd1 vccd1 _09170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08121_ _08323_/A _08323_/B _08120_/X vssd1 vssd1 vccd1 vccd1 _08271_/B sky130_fd_sc_hd__a21o_1
XFILLER_159_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_122_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15464_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08052_ _08052_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08077_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_838 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput109 x_i_6[4] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_1
X_08954_ _15468_/Q _15452_/Q _08953_/X vssd1 vssd1 vccd1 vccd1 _08955_/B sky130_fd_sc_hd__a21oi_2
XFILLER_97_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ _07905_/A vssd1 vssd1 vccd1 vccd1 _15053_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08885_ _15468_/Q _15452_/Q vssd1 vssd1 vccd1 vccd1 _08885_/X sky130_fd_sc_hd__and2b_1
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater840 input65/X vssd1 vssd1 vccd1 vccd1 _07428_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater851 input59/X vssd1 vssd1 vccd1 vccd1 repeater851/X sky130_fd_sc_hd__buf_2
XFILLER_45_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07836_ _15349_/Q input163/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07837_/A sky130_fd_sc_hd__mux2_1
Xrepeater862 input4/X vssd1 vssd1 vccd1 vccd1 _07620_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater873 repeater874/X vssd1 vssd1 vccd1 vccd1 _07663_/A1 sky130_fd_sc_hd__buf_4
Xrepeater884 input240/X vssd1 vssd1 vccd1 vccd1 _07789_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater895 input226/X vssd1 vssd1 vccd1 vccd1 _07720_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07767_ _15383_/Q input155/X _07795_/S vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14169__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _15256_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__08167__A _15012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ _07698_/A vssd1 vssd1 vccd1 vccd1 _15417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _15532_/Q _15516_/Q vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__xnor2_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _15141_/D sky130_fd_sc_hd__xor2_1
XFILLER_40_668 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ _15726_/Q _11431_/B vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__nand2_1
X_09299_ _15403_/Q _15387_/Q vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__xnor2_2
XFILLER_123_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15706_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _14995_/Q vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11261_ _11261_/A _11261_/B vssd1 vssd1 vccd1 vccd1 _11261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14632__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input174_A x_r_2[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _10211_/A _10211_/C _11398_/A vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__a21oi_1
X_13000_ _13273_/A _13201_/A vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11192_ _15750_/Q _15028_/Q vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10143_ _10135_/Y _10139_/B _10137_/B vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__o21ai_1
XFILLER_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A x_i_2[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ _15784_/CLK _14951_/D _13983_/Y vssd1 vssd1 vccd1 vccd1 _14951_/Q sky130_fd_sc_hd__dfrtp_1
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _14982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13902_ _13901_/B _13901_/C _13901_/A vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__o21a_1
X_14882_ _14889_/A vssd1 vssd1 vccd1 vccd1 _14882_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _13832_/A _13832_/C _13832_/B vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14079__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ _13764_/A _13764_/B _13764_/C vssd1 vssd1 vccd1 vccd1 _13765_/B sky130_fd_sc_hd__and3_1
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08077__A _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _15008_/D sky130_fd_sc_hd__nor2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _15572_/CLK _15503_/D _14567_/Y vssd1 vssd1 vccd1 vccd1 _15503_/Q sky130_fd_sc_hd__dfrtp_2
X_12715_ _15052_/Q _12818_/B vssd1 vssd1 vccd1 vccd1 _12827_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ _14976_/Q _13827_/B vssd1 vssd1 vccd1 vccd1 _13696_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14807__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12036__D1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15434_ _15434_/CLK _15434_/D _14494_/Y vssd1 vssd1 vccd1 vccd1 _15434_/Q sky130_fd_sc_hd__dfrtp_2
X_12646_ _12704_/A _12704_/B vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output393_A output393/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15677_/CLK sky130_fd_sc_hd__clkbuf_16
X_15365_ _15374_/CLK _15365_/D _14421_/Y vssd1 vssd1 vccd1 vccd1 _15365_/Q sky130_fd_sc_hd__dfrtp_4
X_12577_ _12575_/A _12575_/B _12576_/X vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__a21oi_2
XFILLER_15_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14316_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14316_/Y sky130_fd_sc_hd__inv_2
X_11528_ _11450_/A _11450_/B _11527_/Y vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__a21oi_1
XFILLER_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15296_ _15563_/CLK _15296_/D _14348_/Y vssd1 vssd1 vccd1 vccd1 _15296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14247_/Y sky130_fd_sc_hd__inv_2
X_11459_ _11537_/B _11459_/B vssd1 vssd1 vccd1 vccd1 _11509_/C sky130_fd_sc_hd__nand2_1
XANTENNA__14542__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater606_A _11363_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14178_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14178_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13712_/A _13712_/B _13713_/B vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__and3_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08670_ _08469_/A _08469_/B _08669_/X vssd1 vssd1 vccd1 vccd1 _08671_/B sky130_fd_sc_hd__o21ai_4
XFILLER_39_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13079__A_N _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A1 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07621_ _07621_/A vssd1 vssd1 vccd1 vccd1 _15455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07552_ _07552_/A vssd1 vssd1 vccd1 vccd1 _15489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07483_ _15522_/Q input23/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07484_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14717__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09222_ _09222_/A _09222_/B _09222_/C vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__and3_1
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09153_ _15564_/Q _15544_/Q vssd1 vssd1 vccd1 vccd1 _09153_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ _11797_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09084_ _09078_/Y _09082_/B _09080_/B vssd1 vssd1 vccd1 vccd1 _09085_/B sky130_fd_sc_hd__o21ai_2
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08035_ _11658_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10695__A_N _15280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput80 x_i_4[7] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
Xinput91 x_i_5[2] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14452__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07765__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _09914_/Y _09985_/B _09916_/B vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__o21ai_1
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ _15462_/Q _15446_/Q vssd1 vssd1 vccd1 vccd1 _08937_/X sky130_fd_sc_hd__and2_1
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08868_ _15466_/Q _15450_/Q vssd1 vssd1 vccd1 vccd1 _08947_/A sky130_fd_sc_hd__xnor2_2
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater670 _14709_/A vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__buf_6
XFILLER_83_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater681 _14515_/A vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_123_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07819_ _07819_/A vssd1 vssd1 vccd1 vccd1 _15358_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater692 _08292_/B vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__buf_6
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ _15342_/Q _15326_/Q vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__nor2_1
XFILLER_189_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10830_ _10828_/A _10828_/B _10829_/X vssd1 vssd1 vccd1 vccd1 _10832_/B sky130_fd_sc_hd__a21o_1
XFILLER_198_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09277__A2 _15381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_900 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12281__A1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ _10768_/A _10761_/B vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__nand2_4
XANTENNA__14627__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_944 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _12500_/A vssd1 vssd1 vccd1 vccd1 _12500_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _10690_/X _10698_/A vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__and2b_2
X_13480_ _13581_/A _13480_/B _13480_/C vssd1 vssd1 vccd1 vccd1 _13481_/B sky130_fd_sc_hd__and3b_1
XFILLER_157_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ _12440_/C _12438_/B _14946_/Q vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15150_ _15394_/CLK _15150_/D _14193_/Y vssd1 vssd1 vccd1 vccd1 _15150_/Q sky130_fd_sc_hd__dfrtp_1
X_12362_ _12371_/A _12371_/C vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__xnor2_2
XFILLER_181_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14101_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__inv_2
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__nor2_2
XFILLER_5_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12293_ _12293_/A vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__clkbuf_2
X_15081_ _15081_/CLK _15081_/D _14121_/Y vssd1 vssd1 vccd1 vccd1 _15081_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14362__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07675__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _11244_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__nand2_1
X_14032_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14032_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08360__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11175_ _11361_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11175_/X sky130_fd_sc_hd__xor2_2
XFILLER_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10126_ _15141_/Q _15306_/Q vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14934_ _15467_/CLK _14934_/D _13965_/Y vssd1 vssd1 vccd1 vccd1 _14934_/Q sky130_fd_sc_hd__dfrtp_1
X_10057_ _15112_/Q _15211_/Q vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__or2b_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14865_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output406_A output406/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11226__A _11226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ _13816_/A _13816_/B vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__and2_1
X_14796_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14796_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12272__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ _13747_/A _13747_/B vssd1 vssd1 vccd1 vccd1 _13748_/C sky130_fd_sc_hd__xnor2_1
XFILLER_56_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10959_ _10959_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _11140_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14537__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater556_A _11289_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ _13672_/A _13672_/B _13677_/X vssd1 vssd1 vccd1 vccd1 _13682_/A sky130_fd_sc_hd__a21oi_2
XFILLER_143_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10784__B _15788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15417_ _15799_/CLK _15417_/D _14476_/Y vssd1 vssd1 vccd1 vccd1 _15417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12629_ _12810_/A _08644_/B _08646_/Y _12628_/Y vssd1 vssd1 vccd1 vccd1 _12648_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _15752_/CLK _15348_/D _14403_/Y vssd1 vssd1 vccd1 vccd1 _15348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07451__A1 _07451_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15279_/CLK _15279_/D _14330_/Y vssd1 vssd1 vccd1 vccd1 _15279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14272__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07585__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _09840_/A _09840_/B _09840_/C vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__and3_1
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09771_/A _09865_/A vssd1 vssd1 vccd1 vccd1 _15725_/D sky130_fd_sc_hd__xnor2_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08653_ _13203_/A _12945_/A vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__xor2_1
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _15463_/Q _07604_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07605_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _08700_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08707_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07535_ _07535_/A vssd1 vssd1 vccd1 vccd1 _15497_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14447__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07466_ _07466_/A vssd1 vssd1 vccd1 vccd1 _15531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _15574_/Q _15554_/Q vssd1 vssd1 vccd1 vccd1 _09205_/Y sky130_fd_sc_hd__nand2_1
XFILLER_210_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07397_ _07397_/A vssd1 vssd1 vccd1 vccd1 _15569_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09136_ _09136_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__or2_1
XFILLER_148_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09067_ _15494_/Q _15478_/Q vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__or2b_1
XFILLER_204_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14182__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08018_ _15800_/Q vssd1 vssd1 vccd1 vccd1 _11898_/A sky130_fd_sc_hd__buf_6
XANTENNA__08180__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09969_ _15201_/Q _15234_/Q vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__xnor2_2
XFILLER_76_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12980_ _15763_/Q _13549_/B vssd1 vssd1 vccd1 vccd1 _13547_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_input137_A x_r_0[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__A_N _15282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11931_/A _11931_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__and3_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14650_/Y sky130_fd_sc_hd__inv_2
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11862_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11866_/C sky130_fd_sc_hd__nor2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _08993_/Y _13600_/B _08995_/B vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__o21ai_2
XFILLER_14_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10813_ _15137_/Q _10812_/Y _10811_/B vssd1 vssd1 vccd1 vccd1 _10814_/B sky130_fd_sc_hd__a21o_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__buf_12
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12403_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14357__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ _12774_/B _13532_/B _13532_/C vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__nand3b_1
X_10744_ _15715_/Q _15781_/Q vssd1 vssd1 vccd1 vccd1 _10744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07681__A1 input182/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13463_ _13463_/A _13463_/B vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__or2_2
X_10675_ _15277_/Q _15178_/Q vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__or2b_1
XANTENNA__08074__B _15792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15202_ _15202_/CLK _15202_/D _14249_/Y vssd1 vssd1 vccd1 vccd1 _15202_/Q sky130_fd_sc_hd__dfrtp_1
X_12414_ _14945_/Q vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__inv_2
XFILLER_142_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _13443_/A _13394_/B vssd1 vssd1 vccd1 vccd1 _13396_/C sky130_fd_sc_hd__or2_1
XFILLER_138_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15133_ _15133_/CLK _15133_/D _14175_/Y vssd1 vssd1 vccd1 vccd1 _15133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12345_ _12246_/B _12330_/S _12130_/B vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09601__B_N _15441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14092__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064_ _15754_/CLK _15064_/D _14103_/Y vssd1 vssd1 vccd1 vccd1 _15064_/Q sky130_fd_sc_hd__dfrtp_1
X_12276_ _12277_/A _12277_/B vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output356_A output356/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14015_/Y sky130_fd_sc_hd__inv_2
X_11227_ _15755_/Q _15033_/Q vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__or2b_1
XFILLER_175_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14820__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _11158_/A _11158_/B vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__nand2_2
XANTENNA_output523_A _15627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ _10109_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_863 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11089_ _14934_/Q _15000_/Q vssd1 vssd1 vccd1 vccd1 _11093_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07434__A _07434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ _15532_/CLK _14917_/D _13947_/Y vssd1 vssd1 vccd1 vccd1 _14917_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14848_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14848_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1052 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12994__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater840_A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15801__D _15801_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14267__A _14269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater938_A input162/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_919 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07424__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14730__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _15089_/Q _15056_/Q vssd1 vssd1 vccd1 vccd1 _09824_/C sky130_fd_sc_hd__or2b_1
XFILLER_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08780__A_N _15337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _09752_/X _09760_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ _13530_/A _08705_/B vssd1 vssd1 vccd1 vccd1 _08706_/A sky130_fd_sc_hd__and2_1
XFILLER_73_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09685_ _09816_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_93_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15750_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08636_ _08711_/A _08588_/Y _08635_/X vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07998__B _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _08567_/A _08629_/B _08567_/C vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__or3_1
XANTENNA__14177__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ _15505_/Q input102/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08498_ _08509_/A _08509_/B vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__xor2_1
XFILLER_195_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07663__A1 _07663_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07449_ _15539_/Q _07449_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07450_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _15159_/Q _15126_/Q vssd1 vssd1 vccd1 vccd1 _10461_/C sky130_fd_sc_hd__or2b_1
XFILLER_13_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _15504_/Q _15488_/Q vssd1 vssd1 vccd1 vccd1 _09258_/A sky130_fd_sc_hd__or2b_1
XFILLER_182_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10391_ _10391_/A _10391_/B _10391_/C vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__and3_1
XANTENNA__12425__A _14945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _12312_/S _12130_/B vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10970__A1 _15269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _12148_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__nand2_1
XFILLER_46_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input254_A x_r_7[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14640__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11012_ _11012_/A _11012_/B vssd1 vssd1 vccd1 vccd1 _15018_/D sky130_fd_sc_hd__xor2_1
XFILLER_81_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15751_ _15752_/CLK _15751_/D _14829_/Y vssd1 vssd1 vccd1 vccd1 _15751_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _13046_/A _12667_/C _12862_/A vssd1 vssd1 vccd1 vccd1 _12963_/X sky130_fd_sc_hd__a21bo_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15712_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__buf_6
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11914_ _12144_/A vssd1 vssd1 vccd1 vccd1 _11991_/A sky130_fd_sc_hd__inv_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15682_ _15687_/CLK _15682_/D _14756_/Y vssd1 vssd1 vccd1 vccd1 _15682_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _13203_/A _12632_/Y _13012_/A vssd1 vssd1 vccd1 vccd1 _12937_/B sky130_fd_sc_hd__mux2_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14633_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14633_/Y sky130_fd_sc_hd__inv_2
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11922_/B _11845_/B vssd1 vssd1 vccd1 vccd1 _11846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14087__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11504__A _15727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14564_/Y sky130_fd_sc_hd__inv_2
X_11776_ _11675_/A _11675_/B _11775_/X vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__a21bo_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12319__B _12323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ _13515_/A _13515_/B vssd1 vssd1 vccd1 vccd1 _15641_/D sky130_fd_sc_hd__xnor2_1
XFILLER_53_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_768 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10727_ _10725_/Y _10727_/B vssd1 vssd1 vccd1 vccd1 _11251_/B sky130_fd_sc_hd__and2b_2
X_14495_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14495_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14815__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13446_ _13463_/B _13446_/B vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__nor2_4
X_10658_ _10652_/A _10654_/B _10652_/B vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__a21boi_4
XANTENNA_output473_A output473/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07406__A1 input124/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13377_ _13438_/A _13390_/A _13491_/S vssd1 vssd1 vccd1 vccd1 _13378_/B sky130_fd_sc_hd__a21o_1
X_10589_ _10589_/A _10628_/A vssd1 vssd1 vccd1 vccd1 _15036_/D sky130_fd_sc_hd__xnor2_1
XFILLER_170_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15116_ _15375_/CLK _15116_/D _14157_/Y vssd1 vssd1 vccd1 vccd1 _15116_/Q sky130_fd_sc_hd__dfrtp_1
X_12328_ _12312_/S _12246_/X _12245_/Y vssd1 vssd1 vccd1 vccd1 _12328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _15493_/CLK _15047_/D _14085_/Y vssd1 vssd1 vccd1 vccd1 _15047_/Q sky130_fd_sc_hd__dfrtp_1
X_12259_ _12207_/Y _12211_/B _12208_/A vssd1 vssd1 vccd1 vccd1 _12260_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14550__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__B1 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater790_A _15602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater888_A repeater889/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12070__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15719_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09470_ _15521_/Q _15537_/Q vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__or2b_1
XFILLER_149_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08421_ _12654_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08426_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ _12357_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__and2_1
XFILLER_177_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08283_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14725__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08723__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12245__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_900 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput530 output530/A vssd1 vssd1 vccd1 vccd1 y_r_7[8] sky130_fd_sc_hd__buf_2
XFILLER_160_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14460__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07773__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _15165_/D sky130_fd_sc_hd__xor2_1
XANTENNA__13076__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07998_ _11797_/A _11658_/A vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_822 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _15064_/Q _15097_/Q vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__xor2_2
XFILLER_39_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09668_ _09667_/A _09667_/C _09667_/B vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08624_/A sky130_fd_sc_hd__and2_1
XANTENNA__07884__A1 input145/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _09597_/X _09604_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__and2b_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11630_ _11630_/A _11697_/C vssd1 vssd1 vccd1 vccd1 _11631_/C sky130_fd_sc_hd__xnor2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07636__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _11618_/B _11561_/B vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14635__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13300_ _13300_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _13301_/B sky130_fd_sc_hd__or2_1
X_10512_ _10512_/A _10512_/B vssd1 vssd1 vccd1 vccd1 _15024_/D sky130_fd_sc_hd__nor2_1
X_14280_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14299_/A sky130_fd_sc_hd__buf_12
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11492_ _11569_/B _11492_/B vssd1 vssd1 vccd1 vccd1 _11493_/C sky130_fd_sc_hd__nand2_1
XFILLER_13_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13231_ _13231_/A _13320_/C vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10443_ _10443_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input65_A x_i_3[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13162_ _13112_/B _13162_/B vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__and2b_1
XFILLER_156_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10374_ _10374_/A _10374_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12113_ _12228_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__or2_1
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14370__A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13203_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07683__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _12160_/A _12044_/B vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__and2_1
XFILLER_105_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _15803_/CLK _15803_/D _14883_/Y vssd1 vssd1 vccd1 vccd1 _15803_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13995_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13995_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15428_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output319_A _15661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ _15790_/CLK _15734_/D _14811_/Y vssd1 vssd1 vccd1 vccd1 _15734_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12946_ _12946_/A _13017_/A vssd1 vssd1 vccd1 vccd1 _13020_/B sky130_fd_sc_hd__xor2_2
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15774_/CLK _15665_/D _14738_/Y vssd1 vssd1 vccd1 vccd1 _15665_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12877_ _12876_/B _12877_/B vssd1 vssd1 vccd1 vccd1 _12878_/B sky130_fd_sc_hd__and2b_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11234__A _15756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14616_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14616_/Y sky130_fd_sc_hd__inv_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11828_/A _11828_/B _11828_/C _11828_/D vssd1 vssd1 vccd1 vccd1 _11829_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_159_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15596_ _15771_/CLK _15596_/D _14666_/Y vssd1 vssd1 vccd1 vccd1 _15596_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14547_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14547_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ _12238_/A _12122_/A vssd1 vssd1 vccd1 vccd1 _12038_/B sky130_fd_sc_hd__xor2_1
XFILLER_186_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14545__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14478_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14478_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13429_ _13380_/A _13380_/B _13385_/A vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__a21o_1
XANTENNA_repeater803_A _15587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _15198_/D sky130_fd_sc_hd__xor2_1
XFILLER_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14280__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07921_ _15429_/Q _15413_/Q vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__or2_1
XFILLER_29_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07852_ _15341_/Q input209/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 enable vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07783_ _15375_/Q _07783_/A1 _07803_/S vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_48_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15663_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09522_ _09522_/A _09522_/B _09522_/C vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__nor3_1
XFILLER_25_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07866__A1 _07866_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _09516_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _15276_/D sky130_fd_sc_hd__xor2_2
XFILLER_149_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09384_ _09382_/X _09386_/C vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__and2b_1
XFILLER_12_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08335_ _11658_/A _11480_/A _08157_/A _11584_/A _08334_/X vssd1 vssd1 vccd1 vccd1
+ _08335_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07618__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14455__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09549__A _15431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08266_ _08279_/A _08279_/B _08265_/X vssd1 vssd1 vccd1 vccd1 _08273_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08453__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08197_ _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14190__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput360 _15684_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[8] sky130_fd_sc_hd__buf_2
XFILLER_134_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput371 _11107_/Y vssd1 vssd1 vccd1 vccd1 y_i_6[2] sky130_fd_sc_hd__buf_2
XFILLER_161_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput382 output382/A vssd1 vssd1 vccd1 vccd1 y_i_7[12] sky130_fd_sc_hd__buf_2
XFILLER_117_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _15215_/Q _15116_/Q _10089_/B vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__a21oi_1
Xoutput393 output393/A vssd1 vssd1 vccd1 vccd1 y_i_7[7] sky130_fd_sc_hd__buf_2
XFILLER_82_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15411_/CLK sky130_fd_sc_hd__clkbuf_16
X_12800_ _12800_/A _12800_/B vssd1 vssd1 vccd1 vccd1 _12800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13780_ _13767_/A _13767_/B _13860_/A _13779_/X vssd1 vssd1 vccd1 vccd1 _13789_/A
+ sky130_fd_sc_hd__o31a_1
X_10992_ _10992_/A _10994_/B vssd1 vssd1 vccd1 vccd1 _15012_/D sky130_fd_sc_hd__nor2_1
XANTENNA_input217_A x_r_5[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _13021_/A vssd1 vssd1 vccd1 vccd1 _12733_/B sky130_fd_sc_hd__inv_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15450_ _15700_/CLK _15450_/D _14511_/Y vssd1 vssd1 vccd1 vccd1 _15450_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__nand2_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14401_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11613_ _11613_/A vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__clkinv_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _15749_/CLK _15381_/D _14437_/Y vssd1 vssd1 vccd1 vccd1 _15381_/Q sky130_fd_sc_hd__dfrtp_4
X_12593_ _12593_/A _12593_/B vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__nand2_1
XFILLER_169_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14365__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14332_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14332_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11544_ _11707_/A _11480_/X _11746_/A _11543_/X vssd1 vssd1 vccd1 vccd1 _11562_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14263_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14263_/Y sky130_fd_sc_hd__inv_2
X_11475_ _11475_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__xnor2_1
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13214_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _15634_/D sky130_fd_sc_hd__nor2_2
XFILLER_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10426_ _10426_/A _10426_/B vssd1 vssd1 vccd1 vccd1 _14950_/D sky130_fd_sc_hd__xor2_2
XFILLER_178_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14194_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14194_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output269_A output269/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__and2_1
X_10357_ _15132_/Q _15165_/Q vssd1 vssd1 vccd1 vccd1 _10359_/A sky130_fd_sc_hd__and2b_1
XFILLER_140_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13352_/A _13366_/A _13076_/C vssd1 vssd1 vccd1 vccd1 _13265_/B sky130_fd_sc_hd__and3_1
XANTENNA__12669__A1 _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__nand2_1
XFILLER_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output436_A _11388_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ _11904_/A _11904_/B _11903_/A _11902_/A _11983_/A vssd1 vssd1 vccd1 vccd1
+ _12126_/B sky130_fd_sc_hd__a311o_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07545__A0 _15492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater586_A repeater587/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _14889_/A vssd1 vssd1 vccd1 vccd1 _13997_/A sky130_fd_sc_hd__buf_12
XFILLER_4_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08538__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15717_ _15717_/CLK _15717_/D _14793_/Y vssd1 vssd1 vccd1 vccd1 _15717_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ _12945_/A _13012_/A vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07848__A1 _07848_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15648_/CLK _15648_/D _14720_/Y vssd1 vssd1 vccd1 vccd1 _15648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15579_ _15680_/CLK _15579_/D _14648_/Y vssd1 vssd1 vccd1 vccd1 _15579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14275__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08120_ _08120_/A _08120_/B _08120_/C vssd1 vssd1 vccd1 vccd1 _08120_/X sky130_fd_sc_hd__and3_1
XFILLER_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08051_ _15802_/Q vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__buf_6
XFILLER_147_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_899 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08953_ _15468_/Q _15452_/Q _08952_/B vssd1 vssd1 vccd1 vccd1 _08953_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07904_ _13874_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07905_/A sky130_fd_sc_hd__and2_1
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07536__A0 _15496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08884_ _08882_/Y _08884_/B vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__nand2b_1
XFILLER_9_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater830 input86/X vssd1 vssd1 vccd1 vccd1 repeater830/X sky130_fd_sc_hd__buf_2
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater841 repeater842/X vssd1 vssd1 vccd1 vccd1 _07430_/A1 sky130_fd_sc_hd__buf_4
X_07835_ _07835_/A vssd1 vssd1 vccd1 vccd1 _15350_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater852 repeater853/X vssd1 vssd1 vccd1 vccd1 _07443_/A1 sky130_fd_sc_hd__buf_4
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater863 input39/X vssd1 vssd1 vccd1 vccd1 _07549_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater874 input254/X vssd1 vssd1 vccd1 vccd1 repeater874/X sky130_fd_sc_hd__buf_2
XFILLER_186_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater885 input24/X vssd1 vssd1 vccd1 vccd1 _07481_/A1 sky130_fd_sc_hd__clkbuf_2
X_07766_ _07766_/A vssd1 vssd1 vccd1 vccd1 _15384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater896 input225/X vssd1 vssd1 vccd1 vccd1 _07722_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08448__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _09421_/Y _09504_/B _09423_/B vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__B _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07697_ _15417_/Q input189/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07698_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09509_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _15273_/D sky130_fd_sc_hd__xor2_1
XFILLER_13_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09365_/A _09365_/B _09366_/X vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14185__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07498__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ _15726_/Q _11431_/B vssd1 vssd1 vccd1 vccd1 _12525_/A sky130_fd_sc_hd__or2_1
XFILLER_177_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ _09365_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _15124_/D sky130_fd_sc_hd__xor2_1
XFILLER_21_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08249_ _08254_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__nor2_1
XFILLER_193_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ _11259_/B _11259_/C _11259_/A vssd1 vssd1 vccd1 vccd1 _11261_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10211_ _10211_/A _11398_/A _10211_/C vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__and3_1
XFILLER_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ _15750_/Q _15028_/Q vssd1 vssd1 vccd1 vccd1 _11191_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input167_A x_r_2[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10142_ _10149_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14950_ _15784_/CLK _14950_/D _13982_/Y vssd1 vssd1 vccd1 vccd1 _14950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10073_ _10071_/X _10079_/A vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__and2b_1
XFILLER_153_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11991__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _13901_/A _13901_/B _13901_/C vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__nor3_1
X_14881_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14881_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_A x_i_1[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13832_ _13832_/A _13832_/B _13832_/C vssd1 vssd1 vccd1 vccd1 _13838_/C sky130_fd_sc_hd__and3_1
XFILLER_78_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _13764_/B _13764_/C _13764_/A vssd1 vssd1 vccd1 vccd1 _13772_/B sky130_fd_sc_hd__a21oi_1
X_10975_ _10974_/B _10974_/C _10974_/A vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__a21oi_1
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__xnor2_1
X_15502_ _15506_/CLK _15502_/D _14566_/Y vssd1 vssd1 vccd1 vccd1 _15502_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_203_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13694_ _13694_/A _13694_/B vssd1 vssd1 vccd1 vccd1 _13827_/B sky130_fd_sc_hd__xor2_4
XFILLER_206_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _15433_/CLK _15433_/D _14493_/Y vssd1 vssd1 vccd1 vccd1 _15433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ _08657_/A _08657_/B _12644_/Y vssd1 vssd1 vccd1 vccd1 _12704_/B sky130_fd_sc_hd__a21o_1
XFILLER_188_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14095__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _15364_/CLK _15364_/D _14419_/Y vssd1 vssd1 vccd1 vccd1 _15364_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_196_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12576_ _14939_/Q _12576_/B vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__and2_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output386_A output386/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14315_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14315_/Y sky130_fd_sc_hd__inv_2
X_11527_ _11527_/A _11527_/B vssd1 vssd1 vccd1 vccd1 _11527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ _15563_/CLK _15295_/D _14347_/Y vssd1 vssd1 vccd1 vccd1 _15295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14246_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14246_/Y sky130_fd_sc_hd__inv_2
X_11458_ _11458_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11459_/B sky130_fd_sc_hd__or2_1
XANTENNA__12354__A3 _08347_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ _10408_/B _10408_/C _10408_/A vssd1 vssd1 vccd1 vccd1 _10412_/B sky130_fd_sc_hd__a21oi_1
X_14177_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14177_/Y sky130_fd_sc_hd__inv_2
X_11389_ _15757_/Q _15035_/Q vssd1 vssd1 vccd1 vccd1 _11389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13128_/A _13128_/B vssd1 vssd1 vccd1 vccd1 _13713_/B sky130_fd_sc_hd__xnor2_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13059_/A _13059_/B vssd1 vssd1 vccd1 vccd1 _13062_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07518__A0 _15505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08730__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _15455_/Q _07620_/A1 _07640_/S vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07551_ _15489_/Q _07551_/A1 _07591_/S vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12814__A1 _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07482_ _07482_/A vssd1 vssd1 vccd1 vccd1 _15523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09221_/A vssd1 vssd1 vccd1 vccd1 _15235_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _09152_/A _09631_/B vssd1 vssd1 vccd1 vccd1 _15286_/D sky130_fd_sc_hd__xnor2_1
XFILLER_159_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08103_ _11876_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08797__A2 _08792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _15497_/Q _15481_/Q vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__14733__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08034_ _15803_/Q vssd1 vssd1 vccd1 vccd1 _12122_/A sky130_fd_sc_hd__buf_6
XFILLER_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput70 x_i_4[12] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput81 x_i_4[8] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_2
Xinput92 x_i_5[3] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_51_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09985_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _14929_/D sky130_fd_sc_hd__xnor2_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08936_ _08936_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _15186_/D sky130_fd_sc_hd__xnor2_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__A _15435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _08945_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _15205_/D sky130_fd_sc_hd__xor2_1
XFILLER_184_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_66_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater660 _14762_/X vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__buf_6
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater671 _14681_/A vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__buf_6
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07818_ _15358_/Q input178/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__mux2_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08178__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater682 _14494_/A vssd1 vssd1 vccd1 vccd1 _14500_/A sky130_fd_sc_hd__buf_6
X_08798_ _13893_/A _08798_/B vssd1 vssd1 vccd1 vccd1 _15077_/D sky130_fd_sc_hd__xor2_1
XFILLER_83_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater693 _08118_/A vssd1 vssd1 vccd1 vccd1 _08530_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_123_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07749_ _07749_/A vssd1 vssd1 vccd1 vccd1 _15392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10760_ _15718_/Q _15784_/Q vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _09418_/Y _15511_/Q _09416_/B vssd1 vssd1 vccd1 vccd1 _09420_/B sky130_fd_sc_hd__a21o_1
XFILLER_186_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _10690_/A _10690_/B _11008_/A vssd1 vssd1 vccd1 vccd1 _10698_/A sky130_fd_sc_hd__a21o_1
XFILLER_179_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_124_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _12455_/B _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__nor3_1
XFILLER_157_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _12355_/A _12355_/B _12360_/X vssd1 vssd1 vccd1 vccd1 _12371_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14643__A _14661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14100_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11312_ _11311_/B _11311_/C _11311_/A vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15081_/CLK _15080_/D _14120_/Y vssd1 vssd1 vccd1 vccd1 _15080_/Q sky130_fd_sc_hd__dfrtp_1
X_12292_ _12500_/A _12292_/B vssd1 vssd1 vccd1 vccd1 _12293_/A sky130_fd_sc_hd__or2_1
XFILLER_4_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14031_/Y sky130_fd_sc_hd__inv_2
X_11243_ _11243_/A _11243_/B vssd1 vssd1 vccd1 vccd1 _11243_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_134_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11544__A1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11174_ _15746_/Q _11173_/Y _11169_/B vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _15141_/Q _15306_/Q vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07691__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ _15483_/CLK _14933_/D _13964_/Y vssd1 vssd1 vccd1 vccd1 _14933_/Q sky130_fd_sc_hd__dfrtp_1
X_10056_ _15211_/Q _15112_/Q vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__or2b_1
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13049__A1 _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14864_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14864_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13815_ _13815_/A _13815_/B vssd1 vssd1 vccd1 vccd1 _15663_/D sky130_fd_sc_hd__xnor2_4
XANTENNA_output301_A output301/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10130__B _15307_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14818__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_733 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13722__A _13722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_50_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_766 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ _13677_/A _13677_/B _13677_/C vssd1 vssd1 vccd1 vccd1 _13677_/X sky130_fd_sc_hd__and3_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10889_ _11113_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__xor2_4
XFILLER_188_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater549_A repeater550/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15416_ _15588_/CLK _15416_/D _14475_/Y vssd1 vssd1 vccd1 vccd1 _15416_/Q sky130_fd_sc_hd__dfrtp_4
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15347_ _15347_/CLK _15347_/D _14402_/Y vssd1 vssd1 vccd1 vccd1 _15347_/Q sky130_fd_sc_hd__dfrtp_2
X_12559_ _12556_/A _12556_/B _12556_/C _12558_/X vssd1 vssd1 vccd1 vccd1 _12560_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_repeater716_A _15703_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14553__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07866__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15278_ _15279_/CLK _15278_/D _14329_/Y vssd1 vssd1 vccd1 vccd1 _15278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14229_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14229_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _15069_/Q _15102_/Q vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__xnor2_2
XFILLER_85_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08725_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__and2_1
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08652_ _13012_/A _12921_/A vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07603_ _07603_/A vssd1 vssd1 vccd1 vccd1 _15464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08583_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08584_/B sky130_fd_sc_hd__or2_1
XANTENNA__14728__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07534_ _15497_/Q input109/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08726__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ _15531_/Q _07465_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_764 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09204_ _09204_/A _09674_/A vssd1 vssd1 vccd1 vccd1 _15297_/D sky130_fd_sc_hd__xor2_1
XFILLER_139_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07396_ _15569_/Q _07396_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09135_ _15508_/Q _15492_/Q vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14463__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09066_ _13631_/A _09064_/B _09065_/X vssd1 vssd1 vccd1 vccd1 _15118_/D sky130_fd_sc_hd__a21o_1
XFILLER_194_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08017_ _11876_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08180__B _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09968_ _09966_/A _10006_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__o21a_1
XANTENNA__12711__A _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08919_ _15474_/Q _15458_/Q vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__and2b_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07805__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _09899_/A vssd1 vssd1 vccd1 vccd1 _14959_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _11931_/A _11931_/B _11931_/C vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__a21o_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11863_/B _11753_/B vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14638__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _15090_/D sky130_fd_sc_hd__xor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _15302_/Q vssd1 vssd1 vccd1 vccd1 _10812_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14580_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14580_/Y sky130_fd_sc_hd__inv_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11789_/A _12540_/A _11791_/Y vssd1 vssd1 vccd1 vccd1 _11873_/B sky130_fd_sc_hd__a21o_1
XFILLER_129_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07540__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _13532_/C _13532_/B _12774_/B vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__a21bo_1
X_10743_ _11265_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_201_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13490_/A _13462_/B vssd1 vssd1 vccd1 vccd1 _13464_/A sky130_fd_sc_hd__nor2_2
XFILLER_90_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10674_ _10994_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _15045_/D sky130_fd_sc_hd__xnor2_4
XANTENNA_input95_A x_i_5[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15201_ _15700_/CLK _15201_/D _14248_/Y vssd1 vssd1 vccd1 vccd1 _15201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12413_ _12413_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _12423_/C sky130_fd_sc_hd__nor2_1
XFILLER_173_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13393_ _13393_/A _13393_/B _13393_/C vssd1 vssd1 vccd1 vccd1 _13394_/B sky130_fd_sc_hd__and3_1
XFILLER_194_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14373__A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15132_ _15133_/CLK _15132_/D _14174_/Y vssd1 vssd1 vccd1 vccd1 _15132_/Q sky130_fd_sc_hd__dfrtp_1
X_12344_ _12230_/B _12327_/S _12108_/B vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__o21a_1
XFILLER_153_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15063_ _15081_/CLK _15063_/D _14102_/Y vssd1 vssd1 vccd1 vccd1 _15063_/Q sky130_fd_sc_hd__dfrtp_1
X_12275_ _12275_/A _12275_/B vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__xnor2_1
XFILLER_126_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14014_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ _11226_/A vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output349_A _15689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _15745_/Q _15023_/Q vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_425 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ _10106_/Y _10108_/B vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11088_ _11088_/A vssd1 vssd1 vccd1 vccd1 _11088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ _10033_/A _10035_/B _10033_/B vssd1 vssd1 vccd1 vccd1 _10040_/B sky130_fd_sc_hd__a21boi_1
X_14916_ _15532_/CLK _14916_/D _13946_/Y vssd1 vssd1 vccd1 vccd1 _14916_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14847_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14847_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater666_A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14548__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1064 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14778_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14778_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater833_A input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ _14978_/Q _13836_/B vssd1 vssd1 vccd1 vccd1 _13729_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14283__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07596__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09096__B _15484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_915 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09753_ _09752_/A _09752_/B _09859_/A vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13346__B _13572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__B1 _13713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _11431_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _15054_/Q _15087_/Q vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__or2b_1
XFILLER_55_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _08711_/A _08588_/Y _08591_/X _08634_/X vssd1 vssd1 vccd1 vccd1 _08635_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14458__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08566_/A _08566_/B _08566_/C vssd1 vssd1 vccd1 vccd1 _08567_/C sky130_fd_sc_hd__and3_1
XFILLER_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ _07517_/A vssd1 vssd1 vccd1 vccd1 _15506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ _13390_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08509_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__A1 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07448_ _07448_/A vssd1 vssd1 vccd1 vccd1 _15540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14193__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ input1/X vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__buf_6
XFILLER_149_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12706__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11747__A1 _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _15488_/Q _15504_/Q vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__or2b_1
XFILLER_129_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _15105_/Q _15204_/Q vssd1 vssd1 vccd1 vccd1 _10391_/C sky130_fd_sc_hd__or2b_1
XFILLER_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09049_ _15362_/Q _15378_/Q vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__and2b_1
XFILLER_190_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _11935_/A _11935_/B _11933_/A _11932_/A _12014_/A vssd1 vssd1 vccd1 vccd1
+ _12148_/B sky130_fd_sc_hd__a311o_1
XFILLER_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11011_ _11010_/A _11010_/B _10697_/B vssd1 vssd1 vccd1 vccd1 _11012_/B sky130_fd_sc_hd__a21o_1
XFILLER_150_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input247_A x_r_7[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15750_/CLK _15750_/D _14828_/Y vssd1 vssd1 vccd1 vccd1 _15750_/Q sky130_fd_sc_hd__dfrtp_2
X_12962_ _13042_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _12965_/A sky130_fd_sc_hd__xnor2_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A x_i_0[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _11928_/A _11913_/B _12008_/A vssd1 vssd1 vccd1 vccd1 _11917_/A sky130_fd_sc_hd__and3_1
X_14701_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14701_/Y sky130_fd_sc_hd__inv_2
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15687_/CLK _15681_/D _14755_/Y vssd1 vssd1 vccd1 vccd1 _15681_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _13203_/A _13273_/A _12893_/C vssd1 vssd1 vccd1 vccd1 _12937_/A sky130_fd_sc_hd__and3_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14368__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11913_/B _11623_/C _12008_/A vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__mux2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14632_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14563_/Y sky130_fd_sc_hd__inv_2
X_11775_ _11775_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__or2b_1
XFILLER_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08300__B1 _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _15711_/Q _15777_/Q vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__nand2_1
X_13514_ _13517_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__nand2_1
XFILLER_207_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14494_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14494_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08851__A1 _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output299_A _10952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ _13445_/A _13445_/B vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__and2_1
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10657_ _10655_/Y _10657_/B vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__and2b_2
XFILLER_139_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13376_ _13491_/S _13438_/A vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__nand2_1
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10588_ _15267_/Q _15300_/Q vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__xnor2_2
XFILLER_126_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output466_A output466/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12327_ _12228_/A _12325_/Y _12327_/S vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__mux2_4
XFILLER_154_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _15375_/CLK _15115_/D _14156_/Y vssd1 vssd1 vccd1 vccd1 _15115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14831__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15046_ _15693_/CLK _15046_/D _14084_/Y vssd1 vssd1 vccd1 vccd1 _15046_/Q sky130_fd_sc_hd__dfrtp_1
X_12258_ _12258_/A vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__inv_2
XANTENNA__12163__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11209_ _11209_/A _11209_/B _11372_/B vssd1 vssd1 vccd1 vccd1 _11209_/X sky130_fd_sc_hd__and3_1
XFILLER_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12254_/A _12204_/A _12312_/S vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__a21o_1
XFILLER_150_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater783_A _15609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater950_A input148/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14278__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08420_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__xor2_1
XFILLER_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _14938_/Q _08351_/B vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__or2_1
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08282_ _08105_/A _08105_/B _08329_/A vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12526__A _15727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08723__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput520 output520/A vssd1 vssd1 vccd1 vccd1 y_r_7[14] sky130_fd_sc_hd__buf_2
XANTENNA__14741__A _14741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput531 _15635_/Q vssd1 vssd1 vccd1 vccd1 y_r_7[9] sky130_fd_sc_hd__buf_2
XFILLER_105_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13357__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12261__A _12262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input2_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _09803_/A _09803_/B _09804_/X vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13076__B _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07997_ _15805_/Q vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_75_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07581__A1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09736_ _09733_/A _09848_/A _09733_/B _09735_/X vssd1 vssd1 vccd1 vccd1 _09739_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_28_834 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _09667_/A _09667_/B _09667_/C vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__and3_1
XANTENNA__14188__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08455_/A _08455_/B _08613_/A vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__o21ai_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08186__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _09597_/A _09597_/B _09799_/A vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__a21o_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_358 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ _08553_/B _08549_/B vssd1 vssd1 vccd1 vccd1 _08550_/B sky130_fd_sc_hd__xnor2_2
XFILLER_11_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _11483_/A _11483_/B _11559_/Y vssd1 vssd1 vccd1 vccd1 _11561_/B sky130_fd_sc_hd__a21oi_1
XFILLER_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10511_ _10510_/A _10510_/C _10596_/A vssd1 vssd1 vccd1 vccd1 _10512_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ _11491_/A _11491_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__or2_1
XFILLER_168_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_920 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input197_A x_r_4[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13320_/C sky130_fd_sc_hd__xnor2_1
X_10442_ _10443_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _14891_/D sky130_fd_sc_hd__xor2_1
XFILLER_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ _13221_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ _15167_/Q _15134_/Q vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__and2b_1
XANTENNA__14651__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12112_ _12228_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input58_A x_i_3[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _13005_/A _13005_/B _13091_/X vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__a21bo_1
XFILLER_2_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12043_ _12042_/A _12042_/B _12042_/C vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__o21ai_1
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _15803_/CLK _15802_/D _14882_/Y vssd1 vssd1 vccd1 vccd1 _15802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13994_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15733_ _15784_/CLK _15733_/D _14810_/Y vssd1 vssd1 vccd1 vccd1 _15733_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A _12945_/B vssd1 vssd1 vccd1 vccd1 _13017_/A sky130_fd_sc_hd__xnor2_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14098__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11515__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15664_/CLK _15664_/D _14737_/Y vssd1 vssd1 vccd1 vccd1 _15664_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12876_ _12877_/B _12876_/B vssd1 vssd1 vccd1 vccd1 _12973_/B sky130_fd_sc_hd__and2b_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__B _15034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14615_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14615_/Y sky130_fd_sc_hd__inv_2
X_11827_ _11612_/A _11827_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11828_/D sky130_fd_sc_hd__and3b_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15764_/CLK _15595_/D _14665_/Y vssd1 vssd1 vccd1 vccd1 _15595_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11766_/A _11758_/B _11758_/C vssd1 vssd1 vccd1 vccd1 _11798_/A sky130_fd_sc_hd__or3_1
XFILLER_109_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14546_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14546_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10709_ _15281_/Q _15182_/Q _10708_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__a21oi_4
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11689_ _11638_/A _11638_/B _11688_/Y vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12346__A _12346_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14477_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14477_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater629_A _11031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13428_ _13428_/A _13428_/B vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__xor2_4
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13359_ _13360_/A _13360_/B vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__nor2_1
XFILLER_155_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07874__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15807__D _15807_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ _15429_/Q _15413_/Q vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15029_ _15498_/CLK _15029_/D _14066_/Y vssd1 vssd1 vccd1 vccd1 _15029_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _07851_/A vssd1 vssd1 vccd1 vccd1 _15342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07563__A1 _07563_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 rst vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_07782_ _07782_/A vssd1 vssd1 vccd1 vccd1 _15376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _15535_/Q _15519_/Q vssd1 vssd1 vccd1 vccd1 _09522_/C sky130_fd_sc_hd__and2_1
XANTENNA__07903__A _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _09514_/A _09446_/B _09451_/X vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__a21o_1
XFILLER_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _08404_/A _08404_/B vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09383_ _09382_/B _09382_/C _09382_/A vssd1 vssd1 vccd1 vccd1 _09386_/C sky130_fd_sc_hd__a21o_1
XFILLER_75_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14736__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08334_ _11584_/A _08157_/A _08331_/X _08332_/X _08333_/Y vssd1 vssd1 vccd1 vccd1
+ _08334_/X sky130_fd_sc_hd__o221a_1
XFILLER_177_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08734__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ _08265_/A _08265_/B _08265_/C vssd1 vssd1 vccd1 vccd1 _08265_/X sky130_fd_sc_hd__and3_1
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08453__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08196_ _08196_/A _11466_/A vssd1 vssd1 vccd1 vccd1 _11467_/B sky130_fd_sc_hd__xnor2_2
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14471__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput350 output350/A vssd1 vssd1 vccd1 vccd1 y_i_5[14] sky130_fd_sc_hd__buf_2
XFILLER_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput361 output361/A vssd1 vssd1 vccd1 vccd1 y_i_5[9] sky130_fd_sc_hd__buf_2
Xoutput372 _11109_/Y vssd1 vssd1 vccd1 vccd1 y_i_6[3] sky130_fd_sc_hd__buf_2
XFILLER_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput383 output383/A vssd1 vssd1 vccd1 vccd1 y_i_7[13] sky130_fd_sc_hd__buf_2
XFILLER_133_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput394 output394/A vssd1 vssd1 vccd1 vccd1 y_i_7[8] sky130_fd_sc_hd__buf_2
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _15061_/Q _15094_/Q vssd1 vssd1 vccd1 vccd1 _09719_/Y sky130_fd_sc_hd__nor2_1
X_10991_ _10990_/B _10990_/C _10990_/A vssd1 vssd1 vccd1 vccd1 _10994_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input112_A x_i_6[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12730_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__or2_1
XFILLER_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08347__C _08347_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12661_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 _12690_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14646__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _11612_/A _11827_/B vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__or2b_1
X_14400_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14419_/A sky130_fd_sc_hd__buf_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _14944_/Q _12591_/B _12588_/B _12395_/Y _12396_/A vssd1 vssd1 vccd1 vccd1
+ _12593_/B sky130_fd_sc_hd__a221o_1
X_15380_ _15741_/CLK _15380_/D _14436_/Y vssd1 vssd1 vccd1 vccd1 _15380_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08644__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ _11480_/A _11617_/A _11478_/B _11707_/A _11906_/A vssd1 vssd1 vccd1 vccd1
+ _11543_/X sky130_fd_sc_hd__o2111a_1
X_14331_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14331_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08363__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14262_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14262_/Y sky130_fd_sc_hd__inv_2
X_11474_ _11906_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__xor2_2
XFILLER_184_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13213_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13214_/B sky130_fd_sc_hd__and3_1
XFILLER_171_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ _15212_/Q _10424_/Y _10423_/B vssd1 vssd1 vccd1 vccd1 _10426_/B sky130_fd_sc_hd__a21o_1
X_14193_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14193_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14381__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13144_ _13120_/B _13144_/B vssd1 vssd1 vccd1 vccd1 _13170_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _15131_/Q _15164_/Q vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07793__A1 _07793_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13180_/A _13075_/B vssd1 vssd1 vccd1 vccd1 _13076_/C sky130_fd_sc_hd__and2_1
X_10287_ _10287_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _15773_/D sky130_fd_sc_hd__xnor2_1
X_12026_ _12439_/B _12427_/B vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__nor2_2
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output331_A output331/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A1 _07545_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output429_A output429/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13977_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13977_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15716_ _15717_/CLK _15716_/D _14792_/Y vssd1 vssd1 vccd1 vccd1 _15716_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12928_ _13002_/A _12928_/B vssd1 vssd1 vccd1 vccd1 _12993_/A sky130_fd_sc_hd__or2_1
XFILLER_74_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__B_N _15785_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15647_ _15649_/CLK _15647_/D _14719_/Y vssd1 vssd1 vccd1 vccd1 _15647_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater746_A _15655_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ _13145_/A _13319_/A _12859_/C vssd1 vssd1 vccd1 vccd1 _12862_/A sky130_fd_sc_hd__and3_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14556__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15578_ _15679_/CLK _15578_/D _14647_/Y vssd1 vssd1 vccd1 vccd1 _15578_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14529_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14529_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater913_A input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _08052_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__or2b_1
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14291__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ _08952_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _15192_/D sky130_fd_sc_hd__xnor2_1
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07903_ _15333_/Q _15317_/Q vssd1 vssd1 vccd1 vccd1 _07904_/B sky130_fd_sc_hd__or2_1
XFILLER_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08883_ _15469_/Q _15453_/Q vssd1 vssd1 vccd1 vccd1 _08884_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07536__A1 input108/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater820 input97/X vssd1 vssd1 vccd1 vccd1 _07461_/A1 sky130_fd_sc_hd__clkbuf_2
X_07834_ _15350_/Q _07834_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07835_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater831 input85/X vssd1 vssd1 vccd1 vccd1 _07455_/A1 sky130_fd_sc_hd__clkbuf_2
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13609__A1 _15372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater842 input64/X vssd1 vssd1 vccd1 vccd1 repeater842/X sky130_fd_sc_hd__buf_2
XFILLER_99_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater853 input58/X vssd1 vssd1 vccd1 vccd1 repeater853/X sky130_fd_sc_hd__buf_2
XFILLER_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater864 input38/X vssd1 vssd1 vccd1 vccd1 _07551_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater875 input253/X vssd1 vssd1 vccd1 vccd1 _07665_/A1 sky130_fd_sc_hd__clkbuf_2
X_07765_ _15384_/Q input156/X _07765_/S vssd1 vssd1 vccd1 vccd1 _07766_/A sky130_fd_sc_hd__mux2_1
Xrepeater886 input238/X vssd1 vssd1 vccd1 vccd1 _07793_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater897 repeater898/X vssd1 vssd1 vccd1 vccd1 _07726_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__08448__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11096__A1 _14935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ _09504_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _15255_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07696_ _07696_/A vssd1 vssd1 vccd1 vccd1 _15418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09435_ _09506_/A _09430_/B _09434_/X vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__a21o_1
XFILLER_73_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14466__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07779__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _15402_/Q _15386_/Q vssd1 vssd1 vccd1 vccd1 _09366_/X sky130_fd_sc_hd__and2b_1
XFILLER_75_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08317_ _08347_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__xnor2_2
XFILLER_127_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _15401_/Q _15385_/Q _09296_/X vssd1 vssd1 vccd1 vccd1 _09298_/B sky130_fd_sc_hd__a21oi_1
XFILLER_201_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08248_ _08289_/A _08288_/A vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__or2_1
XFILLER_181_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12348__A1 _12332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08179_ _08177_/Y _08246_/B _11467_/A vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__mux2_1
XFILLER_165_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ _15237_/Q _15072_/Q vssd1 vssd1 vccd1 vccd1 _10211_/C sky130_fd_sc_hd__or2b_1
XFILLER_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11190_ _11365_/A _11190_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07775__A1 input232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ _15144_/Q _15309_/Q vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ _10071_/A _10071_/B _10426_/A vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13900_ _15343_/Q _15327_/Q vssd1 vssd1 vccd1 vccd1 _13901_/C sky130_fd_sc_hd__and2_1
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11991__C _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_940 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13831_ _14977_/Q _13830_/B _13826_/B _13696_/B _13827_/X vssd1 vssd1 vccd1 vccd1
+ _13832_/C sky130_fd_sc_hd__a221o_1
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _10974_/A _10974_/B _10974_/C vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__and3_1
X_13762_ _13769_/A _13769_/B vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__xnor2_1
XFILLER_204_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15501_/CLK _15501_/D _14565_/Y vssd1 vssd1 vccd1 vccd1 _15501_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_189_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12713_ _13203_/A _13273_/A vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__xor2_2
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14376__A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ _13693_/A _13693_/B vssd1 vssd1 vccd1 vccd1 _13694_/B sky130_fd_sc_hd__and2_2
XFILLER_203_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07689__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12036__B1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15432_ _15803_/CLK _15432_/D _14492_/Y vssd1 vssd1 vccd1 vccd1 _15432_/Q sky130_fd_sc_hd__dfrtp_2
X_12644_ _12644_/A _12644_/B vssd1 vssd1 vccd1 vccd1 _12644_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12575_ _12575_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__xor2_4
X_15363_ _15363_/CLK _15363_/D _14418_/Y vssd1 vssd1 vccd1 vccd1 _15363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_873 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07463__A0 _15532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14314_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14314_/Y sky130_fd_sc_hd__inv_2
X_11526_ _11526_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11585_/B sky130_fd_sc_hd__xor2_1
XFILLER_183_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output281_A output281/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15294_ _15563_/CLK _15294_/D _14346_/Y vssd1 vssd1 vccd1 vccd1 _15294_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _11458_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14245_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14245_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_50 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ _10408_/A _10408_/B _10408_/C vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__and3_1
X_14176_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14176_/Y sky130_fd_sc_hd__inv_2
X_11388_ _11388_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11388_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10339_/A _10473_/A vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__nand2_1
X_13127_ _13059_/A _13059_/B _13126_/X vssd1 vssd1 vccd1 vccd1 _13128_/B sky130_fd_sc_hd__o21ai_2
XFILLER_152_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__A2 _15514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13058_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__and2_1
XFILLER_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07518__A1 input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater696_A _08223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12089_/B _12009_/B vssd1 vssd1 vccd1 vccd1 _12009_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07550_ _07550_/A vssd1 vssd1 vccd1 vccd1 _15490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_207_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ _15523_/Q _07481_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14286__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09220_ _09222_/C _09220_/B vssd1 vssd1 vccd1 vccd1 _09221_/A sky130_fd_sc_hd__and2_1
XFILLER_210_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_738 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ _09151_/A _09151_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ _11876_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__and2_1
XFILLER_159_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09082_ _09227_/A _09082_/B vssd1 vssd1 vccd1 vccd1 _15221_/D sky130_fd_sc_hd__xor2_1
XFILLER_175_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ _08040_/B _08040_/A vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__and2b_1
Xinput60 x_i_3[3] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 x_i_4[13] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput82 x_i_4[9] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput93 x_i_5[4] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07757__A1 _07757_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09909_/A _09983_/B _09909_/B vssd1 vssd1 vccd1 vccd1 _09985_/B sky130_fd_sc_hd__a21boi_1
XFILLER_131_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _08976_/A _08933_/B _08934_/X vssd1 vssd1 vccd1 vccd1 _15217_/D sky130_fd_sc_hd__a21o_1
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13365__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__B _15419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08866_ _08942_/A _08861_/B _08865_/X vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__a21o_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater650 _07971_/Y vssd1 vssd1 vccd1 vccd1 output396/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ _07817_/A vssd1 vssd1 vccd1 vccd1 _15359_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater661 _14781_/A vssd1 vssd1 vccd1 vccd1 _14780_/A sky130_fd_sc_hd__buf_6
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater672 _14675_/A vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__buf_6
X_08797_ _13890_/A _08792_/B _08796_/X vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__a21o_1
XFILLER_177_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater683 _14488_/A vssd1 vssd1 vccd1 vccd1 _14494_/A sky130_fd_sc_hd__buf_6
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08178__B _08223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater694 _14881_/A vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__buf_6
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07748_ _15392_/Q _07748_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07679_ _15426_/Q input183/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14196__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15730__D _15730_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07693__A0 _15419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11097__A_N _14936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _15527_/Q vssd1 vssd1 vccd1 vccd1 _09418_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10690_ _10690_/A _10690_/B _11008_/A vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__and3_1
XFILLER_185_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12342__A_N _12339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _15381_/Q vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__inv_2
XFILLER_200_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07445__A0 _15541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ _11507_/B _12360_/B vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__and2b_1
XFILLER_205_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11311_ _11311_/A _11311_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__and3_1
X_12291_ _12291_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12292_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14030_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14030_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11242_ _11244_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11243_/B sky130_fd_sc_hd__and2_1
XFILLER_84_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07748__A1 _07748_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ _15024_/Q vssd1 vssd1 vccd1 vccd1 _11173_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10124_ _10821_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _15797_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_input40_A x_i_2[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14932_ _15500_/CLK _14932_/D _13963_/Y vssd1 vssd1 vccd1 vccd1 _14932_/Q sky130_fd_sc_hd__dfrtp_1
X_10055_ _10412_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _14979_/D sky130_fd_sc_hd__xnor2_2
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14863_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14863_/Y sky130_fd_sc_hd__inv_2
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_910 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _13812_/A _13812_/B _13813_/X vssd1 vssd1 vccd1 vccd1 _13815_/B sky130_fd_sc_hd__o21ai_2
XFILLER_1_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14794_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14794_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ _13740_/B _13740_/C _13740_/A vssd1 vssd1 vccd1 vccd1 _13748_/B sky130_fd_sc_hd__a21o_1
XFILLER_189_745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ _10959_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__and2_1
XFILLER_43_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_784 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _13674_/A _13819_/A _13675_/X vssd1 vssd1 vccd1 vccd1 _13684_/A sky130_fd_sc_hd__a21o_1
X_10888_ _14958_/Q _10887_/Y _10883_/B vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12338__B _12339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output496_A output496/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15415_ _15799_/CLK _15415_/D _14474_/Y vssd1 vssd1 vccd1 vccd1 _15415_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12627_ _12627_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14834__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15346_ _15346_/CLK _15346_/D _14401_/Y vssd1 vssd1 vccd1 vccd1 _15346_/Q sky130_fd_sc_hd__dfrtp_1
X_12558_ _12154_/B _15736_/Q vssd1 vssd1 vccd1 vccd1 _12558_/X sky130_fd_sc_hd__and2b_1
XFILLER_8_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11509_ _11509_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__nand3_2
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater611_A repeater612/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15277_ _15433_/CLK _15277_/D _14328_/Y vssd1 vssd1 vccd1 vccd1 _15277_/Q sky130_fd_sc_hd__dfrtp_1
X_12489_ _12498_/B _12489_/B vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__and2_1
XFILLER_156_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater709_A _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14228_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14176_/A sky130_fd_sc_hd__buf_6
XFILLER_98_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07882__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater980_A repeater981/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__A2 _13563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08720_ _08715_/Y _08718_/X _08714_/X vssd1 vssd1 vccd1 vccd1 _08720_/X sky130_fd_sc_hd__o21a_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08651_ _15050_/Q vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__buf_4
XFILLER_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07602_ _15464_/Q input76/X _07644_/S vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__mux2_1
XFILLER_208_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08582_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__nand2_2
XFILLER_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _07533_/A vssd1 vssd1 vccd1 vccd1 _15498_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07911__A _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08726__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07464_ _07464_/A vssd1 vssd1 vccd1 vccd1 _15532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09203_ _15574_/Q _15554_/Q vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07395_ _07395_/A vssd1 vssd1 vccd1 vccd1 _15570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14744__A _14751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09134_ _15508_/Q _15492_/Q vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__and2_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _15380_/Q _15364_/Q vssd1 vssd1 vccd1 vccd1 _09065_/X sky130_fd_sc_hd__and2b_1
XFILLER_175_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08016_ _15806_/Q vssd1 vssd1 vccd1 vccd1 _12308_/S sky130_fd_sc_hd__buf_4
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13079__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09573__A _15437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15725__D _15725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _15458_/Q _15474_/Q vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__and2b_1
XFILLER_170_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09904_/A vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__and2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _15446_/Q _15462_/Q vssd1 vssd1 vccd1 vccd1 _08850_/B sky130_fd_sc_hd__and2b_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11935_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__nand2_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10811_/A _10811_/B vssd1 vssd1 vccd1 vccd1 _14906_/D sky130_fd_sc_hd__nor2_1
X_11791_ _11791_/A _12541_/B vssd1 vssd1 vccd1 vccd1 _11791_/Y sky130_fd_sc_hd__nor2_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _13530_/A _13528_/B vssd1 vssd1 vccd1 vccd1 _13532_/B sky130_fd_sc_hd__or2b_1
X_10742_ _10734_/Y _10738_/B _10736_/B vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__o21ai_4
XFILLER_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10673_ _10665_/Y _10669_/B _10667_/B vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__o21ai_4
XFILLER_139_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13461_ _13461_/A _13461_/B _13461_/C vssd1 vssd1 vccd1 vccd1 _13462_/B sky130_fd_sc_hd__and3_1
XFILLER_159_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14654__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ _15763_/CLK _15200_/D _14247_/Y vssd1 vssd1 vccd1 vccd1 _15200_/Q sky130_fd_sc_hd__dfrtp_1
X_12412_ _14944_/Q vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__inv_2
XFILLER_51_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input88_A x_i_5[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08652__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ _13393_/A _13393_/B _13393_/C vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__a21oi_1
X_15131_ _15729_/CLK _15131_/D _14173_/Y vssd1 vssd1 vccd1 vccd1 _15131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12343_ _12341_/A _12571_/A _12342_/X vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12274_ _12308_/S _12230_/X _12231_/B vssd1 vssd1 vccd1 vccd1 _12275_/B sky130_fd_sc_hd__o21ai_1
X_15062_ _15081_/CLK _15062_/D _14101_/Y vssd1 vssd1 vccd1 vccd1 _15062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14013_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14013_/Y sky130_fd_sc_hd__inv_2
X_11225_ _11223_/X _11230_/B vssd1 vssd1 vccd1 vccd1 _11226_/A sky130_fd_sc_hd__and2b_1
XFILLER_136_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11156_ _15745_/Q _15023_/Q vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__or2_1
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ _15137_/Q _15302_/Q vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _11085_/X _11093_/A vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__and2b_1
Xinput250 x_r_7[1] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_1
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ _10036_/Y _10038_/B vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__and2b_1
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14915_ _15532_/CLK _14915_/D _13945_/Y vssd1 vssd1 vccd1 vccd1 _14915_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output411_A output411/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output509_A output509/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14829__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14846_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14777_ _14781_/A vssd1 vssd1 vccd1 vccd1 _14777_/Y sky130_fd_sc_hd__inv_2
X_11989_ _12254_/A _12247_/A _11987_/X vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__a21o_1
XFILLER_17_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07657__A0 _15437_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13728_ _13728_/A _13732_/C vssd1 vssd1 vccd1 vccd1 _13838_/B sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_50_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__B _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13816_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_repeater826_A input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14564__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ _15345_/CLK _15329_/D _14383_/Y vssd1 vssd1 vccd1 vccd1 _15329_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_65_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09821_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _15745_/D sky130_fd_sc_hd__xor2_2
XFILLER_8_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07906__A _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ _09752_/A _09752_/B _09859_/A vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_123_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08703_ _11431_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__or2_1
X_09683_ _15087_/Q _15054_/Q vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__or2b_1
XANTENNA__12958__S _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14739__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _08713_/A _08713_/B _08632_/Y _08633_/Y vssd1 vssd1 vccd1 vccd1 _08634_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08565_ _08629_/A vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15280__D _15280_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07516_ _15506_/Q _07516_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _08496_/A _08520_/C vssd1 vssd1 vccd1 vccd1 _08511_/B sky130_fd_sc_hd__xnor2_1
XFILLER_165_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10998__B_N _15276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11995__A2 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07447_ _15540_/Q _07447_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14474__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08860__A2 _15447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07787__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__A _15436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09117_ _15503_/Q _15487_/Q _09116_/B vssd1 vssd1 vccd1 vccd1 _09121_/A sky130_fd_sc_hd__a21o_1
XFILLER_202_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09048_ _09048_/A vssd1 vssd1 vccd1 vccd1 _15114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ _11010_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _15017_/D sky130_fd_sc_hd__xor2_1
XFILLER_145_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11338__A _11338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input142_A x_r_0[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12961_ _13025_/A _13025_/B vssd1 vssd1 vccd1 vccd1 _13042_/B sky130_fd_sc_hd__xnor2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14649__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11912_ _11912_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11986_/A sky130_fd_sc_hd__xnor2_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15680_ _15680_/CLK _15680_/D _14754_/Y vssd1 vssd1 vccd1 vccd1 _15680_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _13012_/A _12892_/B vssd1 vssd1 vccd1 vccd1 _12896_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1026 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14631_/Y sky130_fd_sc_hd__inv_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _12088_/A vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__inv_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14562_/Y sky130_fd_sc_hd__inv_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11817_/B _11774_/B vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__nand2_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__A1 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__B2 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13513_/A _15772_/Q vssd1 vssd1 vccd1 vccd1 _13517_/A sky130_fd_sc_hd__or2b_1
XFILLER_41_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10725_ _15711_/Q _15777_/Q vssd1 vssd1 vccd1 vccd1 _10725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14493_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14384__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07697__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11801__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13444_ _13445_/A _13445_/B vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ _15273_/Q _15174_/Q vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08382__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1092 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13375_ _13375_/A _13332_/A vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__or2b_1
X_10587_ _10585_/A _10625_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__o21a_1
X_15114_ _15375_/CLK _15114_/D _14155_/Y vssd1 vssd1 vccd1 vccd1 _15114_/Q sky130_fd_sc_hd__dfrtp_1
X_12326_ _12326_/A _12309_/B vssd1 vssd1 vccd1 vccd1 _12327_/S sky130_fd_sc_hd__or2b_1
XFILLER_126_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output361_A output361/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output459_A _15599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ _15508_/CLK _15045_/D _14083_/Y vssd1 vssd1 vccd1 vccd1 _15045_/Q sky130_fd_sc_hd__dfrtp_1
X_12257_ _12257_/A _12257_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__or2_1
XFILLER_170_979 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12632__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12163__A2 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11208_/A _11216_/A vssd1 vssd1 vccd1 vccd1 _11372_/B sky130_fd_sc_hd__nand2_1
X_12188_ _12312_/S _12254_/A vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13447__B _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11139_ _11137_/A _11137_/B _11138_/X vssd1 vssd1 vccd1 vccd1 _11140_/B sky130_fd_sc_hd__a21oi_2
XFILLER_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14559__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater776_A repeater777/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14829_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14829_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater943_A input158/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08350_ _14938_/Q _08351_/B vssd1 vssd1 vccd1 vccd1 _12357_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08281_ _08281_/A _08281_/B vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14294__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08292__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07400__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__A _15127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput510 output510/A vssd1 vssd1 vccd1 vccd1 y_r_6[5] sky130_fd_sc_hd__buf_2
XFILLER_69_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput521 output521/A vssd1 vssd1 vccd1 vccd1 y_r_7[15] sky130_fd_sc_hd__buf_2
XFILLER_172_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13357__B _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15275__D _15275_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09804_ _15441_/Q _15425_/Q vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__and2_1
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07996_ _12178_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08004_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09735_ _15063_/Q _15096_/Q vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__and2_1
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14469__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09666_ _09666_/A vssd1 vssd1 vccd1 vccd1 _15311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _12708_/A _12871_/A _08609_/Y _08611_/X _08616_/Y vssd1 vssd1 vccd1 vccd1
+ _08617_/X sky130_fd_sc_hd__o221a_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09597_/B _09799_/A vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__and3_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08548_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__xnor2_2
XFILLER_126_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08479_ _13319_/A _08531_/B vssd1 vssd1 vccd1 vccd1 _08486_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _10510_/A _10596_/A _10510_/C vssd1 vssd1 vccd1 vccd1 _10512_/A sky130_fd_sc_hd__and3_1
X_11490_ _11491_/A _11491_/B vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _15121_/Q _10440_/Y _10439_/B vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _15134_/Q _15167_/Q vssd1 vssd1 vccd1 vccd1 _10374_/A sky130_fd_sc_hd__and2b_1
XFILLER_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13160_ _13233_/A _13160_/B vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__or2_1
XFILLER_200_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ _12111_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__xor2_1
X_13091_ _13091_/A _13007_/B vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__or2b_1
XFILLER_46_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12042_/A _12042_/B _12042_/C vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__or3_1
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15801_ _15808_/CLK _15801_/D _14881_/Y vssd1 vssd1 vccd1 vccd1 _15801_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13993_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14379__A _14379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ _15732_/CLK _15732_/D _14809_/Y vssd1 vssd1 vccd1 vccd1 _15732_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12942_/Y _12944_/B vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__and2b_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08377__A _15048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15663_ _15663_/CLK _15663_/D _14736_/Y vssd1 vssd1 vccd1 vccd1 _15663_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ _13056_/B _12809_/B _12804_/Y vssd1 vssd1 vccd1 vccd1 _12876_/B sky130_fd_sc_hd__a21o_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14614_/Y sky130_fd_sc_hd__inv_2
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11681_/A _11823_/X _11828_/C _11683_/X _11825_/X vssd1 vssd1 vccd1 vccd1
+ _11829_/B sky130_fd_sc_hd__a221oi_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15761_/CLK _15594_/D _14664_/Y vssd1 vssd1 vccd1 vccd1 _15594_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14545_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ _11678_/A _11678_/B _11756_/Y vssd1 vssd1 vccd1 vccd1 _11825_/B sky130_fd_sc_hd__a21bo_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12627__A _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _15050_/D sky130_fd_sc_hd__nor2_2
XFILLER_119_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_898 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14476_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14476_/Y sky130_fd_sc_hd__inv_2
X_11688_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11688_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ _13370_/B _13372_/B _13370_/A vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__o21ba_2
X_10639_ _10639_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _15038_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__14842__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13422_/A _13357_/Y _13301_/A _13300_/A _13298_/B vssd1 vssd1 vccd1 vccd1
+ _13360_/B sky130_fd_sc_hd__o32a_1
XANTENNA__08840__A _15348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__B1 _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12309_ _12326_/A _12309_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__xor2_4
X_13289_ _13409_/A _13565_/A _13288_/X vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__o21a_1
XFILLER_46_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15028_ _15498_/CLK _15028_/D _14065_/Y vssd1 vssd1 vccd1 vccd1 _15028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07850_ _15342_/Q _07850_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07890__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07781_ _15376_/Q input229/X _07791_/S vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__mux2_1
Xinput3 x_i_0[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14289__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_632 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09520_ _09520_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _15261_/D sky130_fd_sc_hd__nor2_1
XANTENNA__07903__B _15317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09451_ _15533_/Q _15517_/Q vssd1 vssd1 vccd1 vccd1 _09451_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13921__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ _08728_/B _08434_/B _08435_/A _08401_/Y vssd1 vssd1 vccd1 vccd1 _08405_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _09382_/A _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__and3_1
XFILLER_75_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08333_ _11447_/C _11491_/A vssd1 vssd1 vccd1 vccd1 _08333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_125_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15506_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08734__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11441__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08279_/A _08279_/B _08267_/A vssd1 vssd1 vccd1 vccd1 _08264_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08195_ _08213_/A _08213_/B _08194_/Y vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__a21oi_2
XFILLER_203_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14752__A _14753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput340 output340/A vssd1 vssd1 vccd1 vccd1 y_i_4[5] sky130_fd_sc_hd__buf_2
XFILLER_133_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput351 output351/A vssd1 vssd1 vccd1 vccd1 y_i_5[15] sky130_fd_sc_hd__buf_2
Xoutput362 _15812_/X vssd1 vssd1 vccd1 vccd1 y_i_6[0] sky130_fd_sc_hd__buf_2
XFILLER_10_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput373 output373/A vssd1 vssd1 vccd1 vccd1 y_i_6[4] sky130_fd_sc_hd__buf_2
XFILLER_133_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput384 _15706_/Q vssd1 vssd1 vccd1 vccd1 y_i_7[14] sky130_fd_sc_hd__buf_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput395 output395/A vssd1 vssd1 vccd1 vccd1 y_i_7[9] sky130_fd_sc_hd__buf_2
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07979_ _15798_/Q vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__buf_6
XANTENNA__14199__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15733__D _15733_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09718_ _09838_/A _09718_/B vssd1 vssd1 vccd1 vccd1 _15716_/D sky130_fd_sc_hd__xnor2_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08197__A _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__and3_1
XFILLER_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _15568_/Q _15548_/Q vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__and2b_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input105_A x_i_6[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ _12768_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__xor2_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11611_ _11611_/A _11611_/B _11611_/C vssd1 vssd1 vccd1 vccd1 _11827_/B sky130_fd_sc_hd__nand3_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12591_ _14944_/Q _12591_/B vssd1 vssd1 vccd1 vccd1 _12593_/A sky130_fd_sc_hd__or2_1
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_116_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15763_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14330_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14330_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11542_ _11542_/A _11489_/A vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__or2b_1
XFILLER_156_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07490__A1 _07490_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14261_/Y sky130_fd_sc_hd__inv_2
X_11473_ _11928_/A _11832_/A vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input70_A x_i_4[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _15113_/Q vssd1 vssd1 vccd1 vccd1 _10424_/Y sky130_fd_sc_hd__inv_2
X_14192_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14192_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _13058_/A _13058_/B _13125_/A _13125_/B _13059_/A vssd1 vssd1 vccd1 vccd1
+ _13173_/C sky130_fd_sc_hd__a2111o_1
X_10355_ _10355_/A vssd1 vssd1 vccd1 vccd1 _15787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13074_ _13422_/A _15051_/Q vssd1 vssd1 vccd1 vccd1 _13075_/B sky130_fd_sc_hd__or2_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__and2_1
XFILLER_111_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ _15734_/Q _12025_/B vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12910__A _12910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13976_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15715_ _15782_/CLK _15715_/D _14791_/Y vssd1 vssd1 vccd1 vccd1 _15715_/Q sky130_fd_sc_hd__dfrtp_1
X_12927_ _12927_/A _12927_/B vssd1 vssd1 vccd1 vccd1 _12928_/B sky130_fd_sc_hd__and2_1
XFILLER_74_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14837__A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15646_ _15680_/CLK _15646_/D _14718_/Y vssd1 vssd1 vccd1 vccd1 _15646_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12858_ _13046_/A _12858_/B vssd1 vssd1 vccd1 vccd1 _12863_/A sky130_fd_sc_hd__nor2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _11892_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__xnor2_1
XFILLER_203_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15577_ _15699_/CLK _15577_/D _14646_/Y vssd1 vssd1 vccd1 vccd1 _15577_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_repeater641_A _11302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12789_ _13381_/B _13220_/A vssd1 vssd1 vccd1 vccd1 _12859_/C sky130_fd_sc_hd__xor2_1
XFILLER_187_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14528_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14528_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07481__A1 _07481_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14459_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14459_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater906_A input213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14572__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ _08872_/Y _08950_/B _08874_/B vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__o21ai_1
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07902_ _15333_/Q _15317_/Q vssd1 vssd1 vccd1 vccd1 _13874_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ _15469_/Q _15453_/Q vssd1 vssd1 vccd1 vccd1 _08882_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater810 _15577_/Q vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07914__A _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ _07833_/A vssd1 vssd1 vccd1 vccd1 _15351_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater821 input95/X vssd1 vssd1 vccd1 vccd1 _07465_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater832 repeater833/X vssd1 vssd1 vccd1 vccd1 _07457_/A1 sky130_fd_sc_hd__buf_4
Xrepeater843 input63/X vssd1 vssd1 vccd1 vccd1 _07432_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13609__A2 _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater854 repeater855/X vssd1 vssd1 vccd1 vccd1 _07416_/A1 sky130_fd_sc_hd__buf_4
Xrepeater865 repeater866/X vssd1 vssd1 vccd1 vccd1 _07555_/A1 sky130_fd_sc_hd__buf_4
XFILLER_2_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater876 input251/X vssd1 vssd1 vccd1 vccd1 _07669_/A1 sky130_fd_sc_hd__clkbuf_2
X_07764_ _07764_/A vssd1 vssd1 vccd1 vccd1 _15385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater887 input237/X vssd1 vssd1 vccd1 vccd1 _07795_/A1 sky130_fd_sc_hd__buf_4
Xrepeater898 input223/X vssd1 vssd1 vccd1 vccd1 repeater898/X sky130_fd_sc_hd__buf_2
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ _15528_/Q _15512_/Q _09502_/X vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__A2 _15001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07695_ _15418_/Q _07695_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14747__A _14751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09434_ _15530_/Q _15514_/Q vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__and2b_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09365_/A _09365_/B vssd1 vssd1 vccd1 vccd1 _15140_/D sky130_fd_sc_hd__xor2_1
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _08316_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08317_/B sky130_fd_sc_hd__or2_1
XFILLER_36_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ _15401_/Q _15385_/Q _09292_/B vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ _11906_/A _11467_/A vssd1 vssd1 vccd1 vccd1 _08288_/A sky130_fd_sc_hd__nand2_1
XFILLER_166_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14482__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__S _07795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11214__B_N _15753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ _11491_/A _08223_/B vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__xor2_2
XFILLER_137_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15728__D _15728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ _15144_/Q _15309_/Q vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__or2_1
XFILLER_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _10071_/A _10071_/B _10426_/A vssd1 vssd1 vccd1 vccd1 _10071_/X sky130_fd_sc_hd__and3_1
XFILLER_43_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08760__A_N _15318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _14977_/Q _13830_/B vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__or2_1
XFILLER_210_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input222_A x_r_5[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13747_/A _13748_/A _13747_/B vssd1 vssd1 vccd1 vccd1 _13764_/C sky130_fd_sc_hd__a21o_1
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10973_ _15171_/Q _15270_/Q vssd1 vssd1 vccd1 vccd1 _10974_/C sky130_fd_sc_hd__or2b_1
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14657__A _14661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15500_ _15500_/CLK _15500_/D _14564_/Y vssd1 vssd1 vccd1 vccd1 _15500_/Q sky130_fd_sc_hd__dfrtp_1
X_12712_ _13012_/A _13201_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__nand2_1
XFILLER_204_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13692_ _13681_/A _13677_/X _13690_/X vssd1 vssd1 vccd1 vccd1 _13693_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08655__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15431_ _15438_/CLK _15431_/D _14491_/Y vssd1 vssd1 vccd1 vccd1 _15431_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _12643_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12177__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15362_ _15717_/CLK _15362_/D _14417_/Y vssd1 vssd1 vccd1 vccd1 _15362_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12574_ _14938_/Q _12574_/B _12574_/C vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__or3_4
XFILLER_184_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14313_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__xor2_1
XFILLER_141_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07463__A1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ _15563_/CLK _15293_/D _14345_/Y vssd1 vssd1 vccd1 vccd1 _15293_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14392__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14244_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14244_/Y sky130_fd_sc_hd__inv_2
X_11456_ _11456_/A _11510_/A vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__xnor2_1
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output274_A output274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15638__D _15638_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_62 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ _15109_/Q _15208_/Q vssd1 vssd1 vccd1 vccd1 _10408_/C sky130_fd_sc_hd__or2b_1
X_14175_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14175_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11387_ _11385_/A _11385_/B _11386_/X vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__a21oi_2
XFILLER_180_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _13126_/A _13050_/B vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10338_ _15162_/Q _15129_/Q vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__or2b_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output441_A output441/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A _13057_/B _13057_/C _13057_/D vssd1 vssd1 vccd1 vccd1 _13058_/B
+ sky130_fd_sc_hd__nand4_1
X_10269_ _10267_/X _10274_/B vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12008_ _12008_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__or2_1
XFILLER_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater591_A _11324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater689_A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13959_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13959_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14567__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater856_A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07480_ _07480_/A vssd1 vssd1 vccd1 vccd1 _15524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15629_ _15763_/CLK _15629_/D _14700_/Y vssd1 vssd1 vccd1 vccd1 _15629_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_194_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09150_ _15563_/Q _15543_/Q vssd1 vssd1 vccd1 vccd1 _09151_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08101_ _08101_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__xor2_1
XFILLER_33_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ _09077_/A _09076_/B _09076_/A vssd1 vssd1 vccd1 vccd1 _09082_/B sky130_fd_sc_hd__o21ba_1
XFILLER_174_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12815__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ _11658_/A _11458_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__and3_1
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 x_i_2[9] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 x_i_3[4] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput72 x_i_4[14] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 x_i_5[0] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_4
Xinput94 x_i_5[5] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08954__A1 _15468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09983_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _14928_/D sky130_fd_sc_hd__xnor2_1
XFILLER_170_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08934_ _15476_/Q _15460_/Q vssd1 vssd1 vccd1 vccd1 _08934_/X sky130_fd_sc_hd__and2b_1
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08865_ _15464_/Q _15448_/Q vssd1 vssd1 vccd1 vccd1 _08865_/X sky130_fd_sc_hd__and2b_1
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15283__D _15283_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater640 _15810_/X vssd1 vssd1 vccd1 vccd1 output328/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ _15359_/Q _07816_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__mux2_1
Xrepeater651 repeater653/X vssd1 vssd1 vccd1 vccd1 output430/A sky130_fd_sc_hd__buf_4
XFILLER_85_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater662 _14762_/X vssd1 vssd1 vccd1 vccd1 _14781_/A sky130_fd_sc_hd__buf_4
XFILLER_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08796_ _15340_/Q _15324_/Q vssd1 vssd1 vccd1 vccd1 _08796_/X sky130_fd_sc_hd__and2b_1
Xrepeater673 _14642_/X vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__buf_4
XFILLER_26_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater684 _14435_/A vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__buf_6
Xrepeater695 _14861_/A vssd1 vssd1 vccd1 vccd1 _14853_/A sky130_fd_sc_hd__buf_6
X_07747_ _07747_/A vssd1 vssd1 vccd1 vccd1 _15393_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14477__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13381__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07678_ _07678_/A vssd1 vssd1 vccd1 vccd1 _15427_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09417_ _15528_/Q _15512_/Q vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__xnor2_2
XFILLER_197_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07693__A1 input191/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ _09343_/A _09347_/B _09343_/B vssd1 vssd1 vccd1 vccd1 _15135_/D sky130_fd_sc_hd__o21ba_1
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07445__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _15120_/D sky130_fd_sc_hd__nor2_1
XFILLER_201_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12725__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _14990_/Q _14924_/Q vssd1 vssd1 vccd1 vccd1 _11311_/C sky130_fd_sc_hd__or2b_1
XFILLER_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12290_ _12291_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12500_/A sky130_fd_sc_hd__and2_1
XFILLER_107_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _15035_/Q _15757_/Q vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__or2b_1
XANTENNA_input172_A x_r_2[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ _11172_/A _11172_/B vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__nand2_2
XFILLER_106_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _10115_/Y _10119_/B _10117_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__o21ai_1
XFILLER_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input33_A x_i_1[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _15501_/CLK _14931_/D _13962_/Y vssd1 vssd1 vccd1 vccd1 _14931_/Q sky130_fd_sc_hd__dfrtp_1
X_10054_ _10046_/Y _10050_/B _10048_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__o21ai_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _14862_/A vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__buf_8
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_922 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13813_ _13813_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13813_/X sky130_fd_sc_hd__or2_1
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14793_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14387__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13744_ _13744_/A _13744_/B vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ _14903_/Q _14969_/Q vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__or2b_1
XANTENNA__08385__A _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13675_ _13820_/B _14974_/Q vssd1 vssd1 vccd1 vccd1 _13675_/X sky130_fd_sc_hd__and2b_1
X_10887_ _14892_/Q vssd1 vssd1 vccd1 vccd1 _10887_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15414_ _15799_/CLK _15414_/D _14473_/Y vssd1 vssd1 vccd1 vccd1 _15414_/Q sky130_fd_sc_hd__dfrtp_1
X_12626_ _08702_/A _13636_/A _12625_/X vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__a21oi_1
XFILLER_129_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output391_A output391/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_941 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output489_A _15611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15345_ _15345_/CLK _15345_/D _14399_/Y vssd1 vssd1 vccd1 vccd1 _15345_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12557_ _12557_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _15620_/D sky130_fd_sc_hd__nor2_1
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _11506_/X _11501_/B _11507_/X vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15276_ _15433_/CLK _15276_/D _14327_/Y vssd1 vssd1 vccd1 vccd1 _15276_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _12488_/A _12488_/B _12488_/C _12607_/A vssd1 vssd1 vccd1 vccd1 _12489_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14227_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14227_/Y sky130_fd_sc_hd__inv_2
X_11439_ _15807_/Q vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__buf_4
XANTENNA__14850__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater604_A repeater605/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14158_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13145_/A _13109_/B _13220_/A vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__and3_1
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14089_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater973_A input118/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1023 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _13422_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07601_ _07601_/A vssd1 vssd1 vccd1 vccd1 _15465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08581_ _08586_/A _08586_/B _08579_/X _08580_/X vssd1 vssd1 vccd1 vccd1 _08583_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14297__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07532_ _15498_/Q _07532_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07911__B _15349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07675__A1 _07675_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13430__B_N _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ _15532_/Q input96/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09202_ _09200_/A _09667_/B _09201_/X vssd1 vssd1 vccd1 vccd1 _09204_/A sky130_fd_sc_hd__a21oi_2
XFILLER_195_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07394_ _15570_/Q input130/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07395_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _09133_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _15232_/D sky130_fd_sc_hd__xor2_1
XFILLER_194_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09064_ _13631_/A _09064_/B vssd1 vssd1 vccd1 vccd1 _15117_/D sky130_fd_sc_hd__xnor2_1
XFILLER_191_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08015_ _12238_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14760__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13079__C _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13376__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14910__D _14910_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _14969_/D sky130_fd_sc_hd__xnor2_2
XFILLER_131_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08917_ _08917_/A vssd1 vssd1 vccd1 vccd1 _15213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09896_/A _09896_/C _09979_/A vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__o21ai_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_96_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15354_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _15462_/Q _15446_/Q vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13823__B _13824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _15338_/Q _15322_/Q vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__xnor2_2
XFILLER_166_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15741__D _15741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11624__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ _10809_/A _10809_/C _10809_/B vssd1 vssd1 vccd1 vccd1 _10811_/B sky130_fd_sc_hd__a21oi_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _15731_/Q vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__inv_2
XANTENNA__14000__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12439__B _12439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10741_ _10741_/A _10741_/B vssd1 vssd1 vccd1 vccd1 _11265_/A sky130_fd_sc_hd__nand2_4
XFILLER_14_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13460_ _13461_/A _13461_/B _13461_/C vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__a21oi_2
XFILLER_9_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10672_ _10679_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10994_/A sky130_fd_sc_hd__nand2_2
X_12411_ _12423_/A _12411_/B vssd1 vssd1 vccd1 vccd1 _15649_/D sky130_fd_sc_hd__nor2_1
XFILLER_159_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13391_ _13441_/B _13391_/B vssd1 vssd1 vccd1 vccd1 _13393_/C sky130_fd_sc_hd__nand2_1
XFILLER_167_974 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15184_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08652__B _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15130_ _15180_/CLK _15130_/D _14172_/Y vssd1 vssd1 vccd1 vccd1 _15130_/Q sky130_fd_sc_hd__dfrtp_1
X_12342_ _12339_/B _15741_/Q vssd1 vssd1 vccd1 vccd1 _12342_/X sky130_fd_sc_hd__and2b_1
XFILLER_182_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _15758_/CLK _15061_/D _14100_/Y vssd1 vssd1 vccd1 vccd1 _15061_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12273_ _12164_/A _12229_/Y _12230_/X _12308_/S vssd1 vssd1 vccd1 vccd1 _12275_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14670__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14012_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14012_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11224_ _11223_/A _11223_/B _11379_/A vssd1 vssd1 vccd1 vccd1 _11230_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11155_ _11155_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10106_ _15137_/Q _15302_/Q vssd1 vssd1 vccd1 vccd1 _10106_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11086_ _11085_/A _11085_/B _11346_/A vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__a21o_1
Xinput240 x_r_6[7] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__clkbuf_1
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput251 x_r_7[2] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15367_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10037_ _15207_/Q _15108_/Q vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__nand2_1
X_14914_ _15532_/CLK _14914_/D _13944_/Y vssd1 vssd1 vccd1 vccd1 _14914_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14845_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14845_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output404_A output404/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _14781_/A vssd1 vssd1 vccd1 vccd1 _14776_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11988_ _11988_/A _11987_/X vssd1 vssd1 vccd1 vccd1 _11990_/A sky130_fd_sc_hd__or2b_1
XFILLER_189_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__A _15371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13727_ _14979_/Q _13841_/A _13841_/B vssd1 vssd1 vccd1 vccd1 _13732_/C sky130_fd_sc_hd__or3_1
XFILLER_210_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _10938_/A _10938_/B _11131_/A vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater554_A _11341_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14845__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12068__C _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13658_ _13669_/A _13669_/B vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__xnor2_2
X_12609_ _12607_/A _12607_/B _12608_/X vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__a21oi_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater721_A _15697_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ _13585_/A _13587_/Y _13585_/B _13588_/Y vssd1 vssd1 vccd1 vccd1 _13590_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_repeater819_A input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15527_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ _15768_/CLK _15328_/D _14382_/Y vssd1 vssd1 vccd1 vccd1 _15328_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10964__A1 _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _15527_/CLK _15259_/D _14309_/Y vssd1 vssd1 vccd1 vccd1 _15259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14580__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _15055_/Q _09819_/Y _09818_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__a21o_1
XFILLER_99_766 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07906__B _15445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__A2 _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09751_ _09751_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15725_/CLK sky130_fd_sc_hd__clkbuf_16
X_08702_ _08702_/A _13636_/A vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13924__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09682_ _09680_/A _09680_/B _09681_/X vssd1 vssd1 vccd1 vccd1 _15316_/D sky130_fd_sc_hd__a21o_1
XFILLER_55_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _08633_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _08633_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07896__A1 _07896_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08564_ _08629_/A _08629_/B vssd1 vssd1 vccd1 vccd1 _08564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07515_ _07515_/A vssd1 vssd1 vccd1 vccd1 _15507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_744 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08495_ _12970_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _08520_/C sky130_fd_sc_hd__xor2_2
XANTENNA__14755__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ _07446_/A vssd1 vssd1 vccd1 vccd1 _15541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09568__B _15420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08472__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09116_ _09116_/A _09116_/B vssd1 vssd1 vccd1 vccd1 _15228_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07820__A1 _07820_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09047_ _09045_/X _09052_/B vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__and2b_1
XANTENNA__14490__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15736__D _15736_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _14966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 _15648_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__xnor2_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A x_r_0[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08928__A _15476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _11988_/A _11911_/B vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__and2_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12945_/A _12921_/A vssd1 vssd1 vccd1 vccd1 _12892_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14630_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14630_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11928_/A _11906_/A _11842_/C vssd1 vssd1 vccd1 vccd1 _11846_/A sky130_fd_sc_hd__and3_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1038 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14561_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__buf_12
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__nand2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14665__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__A2 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ _13586_/A vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__inv_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _15710_/Q _15776_/Q _10723_/B vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__a21oi_4
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14492_/Y sky130_fd_sc_hd__inv_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11801__B _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ _13443_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13445_/B sky130_fd_sc_hd__nor2_1
XFILLER_201_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10655_ _15273_/Q _15174_/Q vssd1 vssd1 vccd1 vccd1 _10655_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13374_ _13374_/A _13380_/A _13374_/C vssd1 vssd1 vccd1 vccd1 _13386_/A sky130_fd_sc_hd__or3_1
XFILLER_194_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10586_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15113_ _15375_/CLK _15113_/D _14154_/Y vssd1 vssd1 vccd1 vccd1 _15113_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_103_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ _12308_/S _12230_/X _12229_/Y vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15044_ _15044_/CLK _15044_/D _14082_/Y vssd1 vssd1 vccd1 vccd1 _15044_/Q sky130_fd_sc_hd__dfrtp_1
X_12256_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__and3_1
XFILLER_142_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output354_A output354/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12632__B _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11207_ _15030_/Q _15752_/Q vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__or2b_1
X_12187_ _12187_/A _12139_/A vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__or2b_1
XFILLER_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ _14968_/Q _14902_/Q vssd1 vssd1 vccd1 vccd1 _11138_/X sky130_fd_sc_hd__and2_1
XFILLER_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output521_A output521/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_972 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11069_ _11066_/A _11335_/A _11066_/B _11068_/X vssd1 vssd1 vccd1 vccd1 _11072_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15528_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater671_A _14681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A1 _07878_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater769_A _15629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14828_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14828_/Y sky130_fd_sc_hd__inv_2
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14759_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14759_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14575__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07888__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08280_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08280_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_177_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08292__B _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13919__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput500 _11219_/X vssd1 vssd1 vccd1 vccd1 y_r_6[11] sky130_fd_sc_hd__buf_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12823__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput511 output511/A vssd1 vssd1 vccd1 vccd1 y_r_6[6] sky130_fd_sc_hd__buf_2
Xoutput522 output522/A vssd1 vssd1 vccd1 vccd1 y_r_7[16] sky130_fd_sc_hd__buf_2
XFILLER_132_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10343__A _15129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09803_ _09803_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _15164_/D sky130_fd_sc_hd__xor2_1
XFILLER_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _07995_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09734_ _09848_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _15719_/D sky130_fd_sc_hd__xnor2_1
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _09663_/X _09667_/C vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__and2b_1
XFILLER_131_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _08725_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _08616_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09596_ _09596_/A _09604_/A vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08547_ _08728_/A _08539_/B _08540_/A _08546_/Y vssd1 vssd1 vccd1 vccd1 _08553_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14485__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__A _15438_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08478_ _08478_/A _08478_/B vssd1 vssd1 vccd1 vccd1 _08531_/B sky130_fd_sc_hd__xnor2_1
XFILLER_204_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08483__A _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ _07429_/A vssd1 vssd1 vccd1 vccd1 _15549_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ _15154_/Q vssd1 vssd1 vccd1 vccd1 _10440_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ _15133_/Q _15166_/Q _10370_/B vssd1 vssd1 vccd1 vccd1 _10375_/A sky130_fd_sc_hd__a21oi_1
XFILLER_137_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12178_/A _12109_/Y _12110_/S vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _13197_/B _13090_/B vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ _12041_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _12042_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_input252_A x_r_7[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1048 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15800_ _15808_/CLK _15800_/D _14880_/Y vssd1 vssd1 vccd1 vccd1 _15800_/Q sky130_fd_sc_hd__dfrtp_1
X_13992_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13992_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15731_ _15732_/CLK _15731_/D _14808_/Y vssd1 vssd1 vccd1 vccd1 _15731_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _12943_/A _12943_/B vssd1 vssd1 vccd1 vccd1 _12944_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13283__B _13567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15663_/CLK _15662_/D _14735_/Y vssd1 vssd1 vccd1 vccd1 _15662_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ _12874_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__xor2_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11779_/B _11825_/B vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__and2b_1
X_14613_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14613_/Y sky130_fd_sc_hd__inv_2
X_15593_ _15741_/CLK _15593_/D _14663_/Y vssd1 vssd1 vccd1 vccd1 _15593_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14395__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14544_/Y sky130_fd_sc_hd__inv_2
X_11756_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11756_/Y sky130_fd_sc_hd__nand2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08393__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_79_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ _10706_/A _10706_/B _11012_/A vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__a21oi_2
X_14475_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14475_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11687_ _11687_/A _11687_/B vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__nand2_1
XFILLER_105_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_122_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ _13426_/A _13426_/B vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__nand2_2
X_10638_ _10636_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__and2b_2
XANTENNA_output471_A _11300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13357_ _13366_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13357_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10569_ _15264_/Q _15297_/Q vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__or2b_1
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08840__B _15332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ _12230_/X _12229_/Y _12308_/S vssd1 vssd1 vccd1 vccd1 _12309_/B sky130_fd_sc_hd__mux2_2
XFILLER_5_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13288_ _13211_/A _13563_/B _13565_/A _13287_/X vssd1 vssd1 vccd1 vccd1 _13288_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_137_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15027_ _15027_/CLK _15027_/D _14064_/Y vssd1 vssd1 vccd1 vccd1 _15027_/Q sky130_fd_sc_hd__dfrtp_1
X_12239_ _12240_/A _12240_/B _12240_/C vssd1 vssd1 vccd1 vccd1 _12239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10163__A _10163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13474__A _13781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07780_ _07780_/A vssd1 vssd1 vccd1 vccd1 _15377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08568__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 x_i_0[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09450_ _09450_/A vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ _08401_/A _08437_/A vssd1 vssd1 vccd1 vccd1 _08401_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ _15406_/Q _15390_/Q vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__or2b_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12818__A _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08332_ _11458_/A _08177_/Y _08330_/Y _11435_/A vssd1 vssd1 vccd1 vccd1 _08332_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12072__A2 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11441__B _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _08194_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _08194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09776__A1 _15431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07787__A0 _15373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput330 output330/A vssd1 vssd1 vccd1 vccd1 y_i_4[11] sky130_fd_sc_hd__buf_2
Xoutput341 output341/A vssd1 vssd1 vccd1 vccd1 y_i_4[6] sky130_fd_sc_hd__buf_2
XFILLER_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput352 output352/A vssd1 vssd1 vccd1 vccd1 y_i_5[16] sky130_fd_sc_hd__buf_2
Xoutput363 output363/A vssd1 vssd1 vccd1 vccd1 y_i_6[10] sky130_fd_sc_hd__buf_2
XFILLER_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput374 output374/A vssd1 vssd1 vccd1 vccd1 y_i_6[5] sky130_fd_sc_hd__buf_2
XFILLER_0_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput385 output385/A vssd1 vssd1 vccd1 vccd1 y_i_7[15] sky130_fd_sc_hd__buf_2
XFILLER_142_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput396 output396/A vssd1 vssd1 vccd1 vccd1 y_r_0[0] sky130_fd_sc_hd__buf_2
XFILLER_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07978_ _15795_/Q vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _09709_/Y _09713_/B _09711_/B vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__o21ai_1
XFILLER_19_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _15307_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _15438_/Q _15422_/Q vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__and2_1
XFILLER_128_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11610_ _11611_/A _11611_/B _11611_/C vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__a21oi_1
XFILLER_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12590_ _12590_/A _12590_/B vssd1 vssd1 vccd1 vccd1 _15682_/D sky130_fd_sc_hd__xor2_2
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11541_ _11828_/A _11828_/B _11827_/C vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__a21oi_2
XFILLER_129_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14269_/A sky130_fd_sc_hd__buf_6
XFILLER_51_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11472_ _15019_/Q vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__buf_4
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13211_ _13211_/A _13563_/B vssd1 vssd1 vccd1 vccd1 _13213_/C sky130_fd_sc_hd__xnor2_1
X_10423_ _10423_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _14949_/D sky130_fd_sc_hd__nor2_1
X_14191_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14191_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_914 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13142_ _13126_/X _13123_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13173_/B sky130_fd_sc_hd__a21o_1
XANTENNA_input63_A x_i_3[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10354_ _10352_/X _10360_/A vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13073_ _13422_/A _15051_/Q vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10285_ _15249_/Q _15084_/Q vssd1 vssd1 vccd1 vccd1 _10288_/B sky130_fd_sc_hd__or2b_1
XFILLER_152_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12024_ _12024_/A vssd1 vssd1 vccd1 vccd1 _15585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13975_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13975_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output317_A output317/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15714_ _15782_/CLK _15714_/D _14790_/Y vssd1 vssd1 vccd1 vccd1 _15714_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12926_ _12927_/A _12927_/B vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__nor2_1
XFILLER_185_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15645_ _15679_/CLK _15645_/D _14717_/Y vssd1 vssd1 vccd1 vccd1 _15645_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _12970_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__nand2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12638__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08835__B _15331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _11808_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__xor2_1
XFILLER_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15576_ _15576_/CLK _15576_/D _14645_/Y vssd1 vssd1 vccd1 vccd1 _15576_/Q sky130_fd_sc_hd__dfrtp_1
X_12788_ _13145_/A _13319_/A vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__nand2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11739_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11835_/A sky130_fd_sc_hd__inv_2
X_14527_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14527_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater634_A _11253_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14853__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14458_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14458_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _13409_/A _13565_/A _13570_/A _13574_/A vssd1 vssd1 vccd1 vccd1 _13409_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_repeater801_A _15590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14389_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14389_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _15191_/D sky130_fd_sc_hd__xor2_1
XFILLER_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07901_ _07901_/A vssd1 vssd1 vccd1 vccd1 _15317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08881_ _08952_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _15208_/D sky130_fd_sc_hd__xor2_2
Xrepeater800 repeater801/X vssd1 vssd1 vccd1 vccd1 output417/A sky130_fd_sc_hd__buf_4
XFILLER_116_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08733__A2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater811 repeater812/X vssd1 vssd1 vccd1 vccd1 output413/A sky130_fd_sc_hd__buf_4
X_07832_ _15351_/Q input171/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07833_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12312__S _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater822 input94/X vssd1 vssd1 vccd1 vccd1 _07467_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater833 input84/X vssd1 vssd1 vccd1 vccd1 repeater833/X sky130_fd_sc_hd__buf_2
Xrepeater844 repeater845/X vssd1 vssd1 vccd1 vccd1 _07435_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__07406__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater855 input56/X vssd1 vssd1 vccd1 vccd1 repeater855/X sky130_fd_sc_hd__buf_2
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater866 input36/X vssd1 vssd1 vccd1 vccd1 repeater866/X sky130_fd_sc_hd__buf_2
X_07763_ _15385_/Q _07763_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07764_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater877 input25/X vssd1 vssd1 vccd1 vccd1 _07479_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_452 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater888 repeater889/X vssd1 vssd1 vccd1 vccd1 _07799_/A1 sky130_fd_sc_hd__buf_4
X_09502_ _15528_/Q _15512_/Q _09501_/B vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13932__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater899 input221/X vssd1 vssd1 vccd1 vccd1 _07730_/A1 sky130_fd_sc_hd__clkbuf_2
X_07694_ _07694_/A vssd1 vssd1 vccd1 vccd1 _15419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07930__A _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ _09431_/Y _09433_/B vssd1 vssd1 vccd1 vccd1 _09509_/A sky130_fd_sc_hd__nand2b_1
XFILLER_198_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ _09362_/A _09362_/B _09363_/X vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ _08322_/A _08275_/B _08313_/Y _08314_/Y vssd1 vssd1 vccd1 vccd1 _08316_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_178_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09295_ _09293_/Y _09295_/B vssd1 vssd1 vccd1 vccd1 _09365_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__14763__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08246_ _11928_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13379__A _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08177_ _11491_/A vssd1 vssd1 vccd1 vccd1 _08177_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__nor2_2
XFILLER_114_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14003__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _13747_/A _13747_/B _13740_/B _13740_/C _13740_/A vssd1 vssd1 vccd1 vccd1
+ _13764_/B sky130_fd_sc_hd__a221o_1
XFILLER_210_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10972_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input215_A x_r_5[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A1 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_934 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _15051_/Q _12711_/B vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13691_ _13681_/A _13690_/X _13672_/A _13672_/B vssd1 vssd1 vccd1 vccd1 _13693_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _15438_/CLK _15430_/D _14490_/Y vssd1 vssd1 vccd1 vccd1 _15430_/Q sky130_fd_sc_hd__dfrtp_1
X_12642_ _12718_/A _12718_/B vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12036__A2 _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15361_ _15719_/CLK _15361_/D _14416_/Y vssd1 vssd1 vccd1 vccd1 _15361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _12573_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _15626_/D sky130_fd_sc_hd__xnor2_1
XFILLER_106_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14673__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11524_ _12228_/A _11600_/B vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14312_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14312_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15292_ _15573_/CLK _15292_/D _14344_/Y vssd1 vssd1 vccd1 vccd1 _15292_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14243_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14243_/Y sky130_fd_sc_hd__inv_2
X_11455_ _08027_/A _08025_/X _08026_/A vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__a21oi_1
XFILLER_7_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10406_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10408_/B sky130_fd_sc_hd__nand2_1
X_14174_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14174_/Y sky130_fd_sc_hd__inv_2
X_11386_ _15756_/Q _15034_/Q vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__and2_1
XFILLER_194_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output267_A _11104_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ _13125_/A _13125_/B vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__nor2_2
X_10337_ _15129_/Q _15162_/Q vssd1 vssd1 vccd1 vccd1 _10339_/A sky130_fd_sc_hd__or2b_1
XFILLER_97_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12921__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13056_ _12804_/Y _13056_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _13057_/D sky130_fd_sc_hd__and3b_1
XANTENNA__13736__B _13746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10268_ _10267_/A _10267_/B _11418_/A vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__a21o_1
XANTENNA_output434_A output434/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_706 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12007_ _12008_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12089_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _15760_/D sky130_fd_sc_hd__nor2_1
XFILLER_120_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11256__B _11257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_867 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater584_A _11125_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14848__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13958_ _14889_/A vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__buf_12
XFILLER_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater751_A repeater752/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _13020_/A _12909_/B _13018_/B vssd1 vssd1 vccd1 vccd1 _12910_/C sky130_fd_sc_hd__nand3_2
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ _08783_/Y _13888_/B _08785_/B vssd1 vssd1 vccd1 vccd1 _13890_/B sky130_fd_sc_hd__o21ai_2
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15628_ _15761_/CLK _15628_/D _14699_/Y vssd1 vssd1 vccd1 vccd1 _15628_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_948 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15559_ _15569_/CLK _15559_/D _14626_/Y vssd1 vssd1 vccd1 vccd1 _15560_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_203_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14583__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _08109_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07896__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _09078_/Y _09080_/B vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__nand2b_2
XFILLER_174_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12815__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08031_ _11678_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__xor2_1
XFILLER_190_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 x_i_2[14] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_880 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput51 x_i_3[0] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput62 x_i_3[5] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput73 x_i_4[15] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
Xinput84 x_i_5[10] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput95 x_i_5[6] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13927__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__A2 _15452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _09900_/Y _09981_/B _09902_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__o21ai_1
XFILLER_116_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08933_ _08976_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _15216_/D sky130_fd_sc_hd__xnor2_1
XFILLER_130_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11447__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08864_ _08862_/Y _08864_/B vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__nand2b_1
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater630 _10875_/X vssd1 vssd1 vccd1 vccd1 output304/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ _07815_/A vssd1 vssd1 vccd1 vccd1 _15360_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater641 _11302_/X vssd1 vssd1 vccd1 vccd1 output336/A sky130_fd_sc_hd__clkbuf_2
Xrepeater652 _07966_/X vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _08793_/Y _08795_/B vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__14758__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater663 _14753_/A vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__buf_6
XFILLER_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07390__A1 _07390_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater674 _14642_/X vssd1 vssd1 vccd1 vccd1 _14661_/A sky130_fd_sc_hd__buf_4
XFILLER_26_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater685 _14439_/A vssd1 vssd1 vccd1 vccd1 _14435_/A sky130_fd_sc_hd__buf_6
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07746_ _15393_/Q _07746_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater696 _08223_/B vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08756__A _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__B _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07677_ _15427_/Q _07677_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08475__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09416_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _15269_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09347_ _09403_/A _09347_/B vssd1 vssd1 vccd1 vccd1 _15134_/D sky130_fd_sc_hd__xor2_4
XFILLER_194_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14493__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11910__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _15397_/Q _15381_/Q _09351_/C vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__and3_1
XANTENNA__08491__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15739__D _15739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ _08292_/B _08236_/B _08237_/A _08228_/Y vssd1 vssd1 vccd1 vccd1 _08232_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _15757_/Q _15035_/Q vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13702__B_N _13062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _15747_/Q _15025_/Q vssd1 vssd1 vccd1 vccd1 _11172_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input165_A x_r_2[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _10122_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__nand2_2
XFILLER_171_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13556__B _13558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14930_ _15501_/CLK _14930_/D _13961_/Y vssd1 vssd1 vccd1 vccd1 _14930_/Q sky130_fd_sc_hd__dfrtp_1
X_10053_ _10060_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__nand2_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A x_i_1[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14861_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14668__A _14681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13572__A _13572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _15662_/D sky130_fd_sc_hd__xor2_4
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14792_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10955_ _14969_/Q _14903_/Q vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__or2b_1
X_13743_ _13743_/A _13842_/A vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__xor2_1
XANTENNA__12188__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _13674_/A _13819_/A vssd1 vssd1 vccd1 vccd1 _15696_/D sky130_fd_sc_hd__xor2_2
XFILLER_204_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15413_ _15803_/CLK _15413_/D _14472_/Y vssd1 vssd1 vccd1 vccd1 _15413_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _13634_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__and2b_1
XFILLER_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12556_ _12556_/A _12556_/B _12556_/C vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__and3_1
XFILLER_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15344_ _15768_/CLK _15344_/D _14398_/Y vssd1 vssd1 vccd1 vccd1 _15344_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output384_A _15706_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _12360_/B _11507_/B vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__and2_1
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12487_ _12488_/A _12488_/B _12488_/C _12607_/A vssd1 vssd1 vccd1 vccd1 _12498_/B
+ sky130_fd_sc_hd__a31o_1
X_15275_ _15433_/CLK _15275_/D _14326_/Y vssd1 vssd1 vccd1 vccd1 _15275_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11438_ _12308_/S _11438_/B vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__nand2_1
X_14226_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14226_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14157_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11369_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13108_ _13235_/B _13108_/B vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__nor2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13040_/A _13040_/B vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10171__A _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater966_A input125/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14578__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07600_ _15465_/Q _07600_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08580_ _08556_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08580_/X sky130_fd_sc_hd__and2b_1
XFILLER_93_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_580 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07531_ _07531_/A vssd1 vssd1 vccd1 vccd1 _15499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_915 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ _07462_/A vssd1 vssd1 vccd1 vccd1 _15533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09201_ _15573_/Q _15553_/Q vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__and2_1
X_07393_ _07393_/A vssd1 vssd1 vccd1 vccd1 _15571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09132_ _15507_/Q _15491_/Q vssd1 vssd1 vccd1 vccd1 _09266_/B sky130_fd_sc_hd__xor2_1
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10703__A_N _15281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _09062_/Y _15363_/Q _09058_/B vssd1 vssd1 vccd1 vccd1 _09064_/B sky130_fd_sc_hd__a21oi_1
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__xor2_1
XFILLER_200_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13376__B _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__and2_1
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08916_ _08914_/X _08921_/B vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__and2b_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09896_ _09896_/A _09979_/A _09896_/C vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__or3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _15445_/Q vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__inv_2
XANTENNA__14488__A _14488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _13883_/A _08778_/B vssd1 vssd1 vccd1 vccd1 _15073_/D sky130_fd_sc_hd__xor2_1
XFILLER_205_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _07729_/A vssd1 vssd1 vccd1 vccd1 _15402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _15714_/Q _15780_/Q vssd1 vssd1 vccd1 vccd1 _10741_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10671_ _15276_/Q _15177_/Q vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11640__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _12410_/A _12590_/A _12410_/C vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__nor3_1
XFILLER_159_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _13390_/A _13390_/B vssd1 vssd1 vccd1 vccd1 _13391_/B sky130_fd_sc_hd__or2_1
XFILLER_90_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _12341_/A _12571_/A vssd1 vssd1 vccd1 vccd1 _15592_/D sky130_fd_sc_hd__xor2_4
XFILLER_51_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_945 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15060_ _15345_/CLK _15060_/D _14098_/Y vssd1 vssd1 vccd1 vccd1 _15060_/Q sky130_fd_sc_hd__dfrtp_1
X_12272_ _12238_/A _12238_/B _12237_/A vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__a21o_1
XFILLER_175_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14011_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14011_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _11223_/A _11223_/B _11379_/A vssd1 vssd1 vccd1 vccd1 _11223_/X sky130_fd_sc_hd__and3_1
XFILLER_135_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ _11153_/A _11153_/B _11355_/A vssd1 vssd1 vccd1 vccd1 _11155_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _15136_/Q _15301_/Q _10103_/Y _10104_/Y vssd1 vssd1 vccd1 vccd1 _10109_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11085_ _11085_/A _11085_/B _11346_/A vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__and3_1
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput230 x_r_6[12] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput241 x_r_6[8] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11227__B_N _15033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput252 x_r_7[3] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10036_ _15207_/Q _15108_/Q vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__nor2_1
X_14913_ _15532_/CLK _14913_/D _13943_/Y vssd1 vssd1 vccd1 vccd1 _14913_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14398__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09274__B_N _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_889 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14844_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__A _08396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07504__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14775_ _14781_/A vssd1 vssd1 vccd1 vccd1 _14775_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _12312_/S _12244_/A vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__xor2_1
XFILLER_90_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11989__A1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13841_/A _13841_/B _14979_/Q vssd1 vssd1 vccd1 vccd1 _13728_/A sky130_fd_sc_hd__o21ai_1
X_10938_ _10938_/A _10938_/B _11131_/A vssd1 vssd1 vccd1 vccd1 _10938_/X sky130_fd_sc_hd__and3_1
XFILLER_205_887 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10869_ _10869_/A _10869_/B vssd1 vssd1 vccd1 vccd1 _10869_/Y sky130_fd_sc_hd__nor2_1
X_13657_ _13651_/A _13656_/Y _13651_/B _13648_/A vssd1 vssd1 vccd1 vccd1 _13659_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_158_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ _14950_/Q _12608_/B vssd1 vssd1 vccd1 vccd1 _12608_/X sky130_fd_sc_hd__and2_1
XFILLER_158_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08606__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13588_ _15773_/Q _13588_/B vssd1 vssd1 vccd1 vccd1 _13588_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08606__B2 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ _15768_/CLK _15327_/D _14381_/Y vssd1 vssd1 vccd1 vccd1 _15327_/Q sky130_fd_sc_hd__dfrtp_1
X_12539_ _12536_/A _12537_/A _12536_/B _12538_/X vssd1 vssd1 vccd1 vccd1 _12540_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_repeater714_A _15705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14861__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10964__A2 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15258_ _15527_/CLK _15258_/D _14308_/Y vssd1 vssd1 vccd1 vccd1 _15258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14209_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14209_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _15221_/CLK _15189_/D _14234_/Y vssd1 vssd1 vccd1 vccd1 _15189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_691 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_745 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09750_ _15099_/Q _15066_/Q vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__and2b_1
XFILLER_140_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08701_ _13634_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__xnor2_4
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09681_ _15576_/Q _15556_/Q vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08632_ _08633_/A _08633_/B _08631_/X vssd1 vssd1 vccd1 vccd1 _08632_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14101__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07414__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _08566_/A _08566_/C vssd1 vssd1 vccd1 vccd1 _08629_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09098__A1 _15499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13940__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ _15507_/Q _07514_/A1 _07538_/S vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08494_ _14910_/Q vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__buf_6
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07445_ _15541_/Q input51/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07446_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ _09114_/A _09114_/C _09250_/A vssd1 vssd1 vccd1 vccd1 _09116_/B sky130_fd_sc_hd__o21a_1
XFILLER_182_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_783 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14771__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09046_ _09045_/A _09045_/B _13622_/A vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12291__A _12291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09948_ _09946_/X _09953_/B vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__and2b_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _15188_/Q _15221_/Q vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _12254_/A _12247_/A vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__or2_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input128_A x_i_7[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12930_/B _12923_/B vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14011__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _12002_/B _11841_/B vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__nor2_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__A1 _15497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__or2_1
XFILLER_14_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14560_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14560_/Y sky130_fd_sc_hd__inv_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10723_ _10723_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10723_/Y sky130_fd_sc_hd__nor2_2
XFILLER_13_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13511_ _15773_/Q _13588_/B vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14491_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14491_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12466__A _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ _10980_/A _10654_/B vssd1 vssd1 vccd1 vccd1 _15041_/D sky130_fd_sc_hd__xnor2_4
XFILLER_139_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13442_ _13463_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__or2_1
XANTENNA_input93_A x_i_5[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ _13373_/A _13343_/B vssd1 vssd1 vccd1 vccd1 _13396_/B sky130_fd_sc_hd__or2b_1
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10585_ _10585_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _15035_/D sky130_fd_sc_hd__xnor2_1
XFILLER_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14681__A _14681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _15363_/CLK _15112_/D _14153_/Y vssd1 vssd1 vccd1 vccd1 _15112_/Q sky130_fd_sc_hd__dfrtp_1
X_12324_ _12321_/A _12322_/X _12323_/X vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__a21o_2
XFILLER_155_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12255_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__a21oi_1
XFILLER_182_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15043_ _15467_/CLK _15043_/D _14081_/Y vssd1 vssd1 vccd1 vccd1 _15043_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10714__A _15282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ _15752_/Q _15030_/Q vssd1 vssd1 vccd1 vccd1 _11208_/A sky130_fd_sc_hd__or2b_1
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12186_ _12186_/A _12137_/B vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__or2b_1
XANTENNA_output347_A _15687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07575__A1 _07575_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ _11137_/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__xor2_4
XFILLER_205_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11068_ _14931_/Q _14997_/Q vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__and2_1
XANTENNA_output514_A _11203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15662__D _15662_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10019_ _10017_/Y _10019_/B vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__and2b_1
XFILLER_209_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14827_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14827_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14856__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater664_A _14750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14758_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08854__A _15463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _13706_/A _13829_/A _13708_/Y vssd1 vssd1 vccd1 vccd1 _13721_/A sky130_fd_sc_hd__a21oi_2
XFILLER_204_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater831_A input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14689_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14689_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater929_A input176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_794 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14591__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput501 _11226_/X vssd1 vssd1 vccd1 vccd1 y_r_6[12] sky130_fd_sc_hd__buf_2
Xoutput512 _11189_/X vssd1 vssd1 vccd1 vccd1 y_r_6[7] sky130_fd_sc_hd__buf_2
XFILLER_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput523 _15627_/Q vssd1 vssd1 vccd1 vccd1 y_r_7[1] sky130_fd_sc_hd__buf_2
XANTENNA__07917__B _15509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13887__A1 _15338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13000__A _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09802_ _15440_/Q _15424_/Q _09801_/B vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13935__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07994_ _11678_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _07995_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ _09663_/A _09663_/C _09663_/B vssd1 vssd1 vccd1 vccd1 _09667_/C sky130_fd_sc_hd__a21o_1
XFILLER_28_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08615_ _08615_/A _08615_/B vssd1 vssd1 vccd1 vccd1 _08721_/B sky130_fd_sc_hd__nand2_1
X_09595_ _15440_/Q _15424_/Q vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__or2b_1
XANTENNA__14766__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08477_ _14914_/Q vssd1 vssd1 vccd1 vccd1 _13319_/A sky130_fd_sc_hd__buf_6
XANTENNA__14916__D _14916_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08483__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07428_ _15549_/Q _07428_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09444__A_N _15532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10370_ _10370_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _15789_/D sky130_fd_sc_hd__nor2_1
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15747__D _15747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09029_ _15375_/Q _15359_/Q vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__or2b_1
XFILLER_151_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14006__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ _12040_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07557__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13845__A _13845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input245_A x_r_7[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13991_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13991_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15730_ _15732_/CLK _15730_/D _14807_/Y vssd1 vssd1 vccd1 vccd1 _15730_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12942_ _12943_/A _12943_/B vssd1 vssd1 vccd1 vccd1 _12942_/Y sky130_fd_sc_hd__nor2_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15677_/CLK _15661_/D _14734_/Y vssd1 vssd1 vccd1 vccd1 _15661_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12873_ _12803_/A _12803_/B _12872_/X vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__a21bo_1
XFILLER_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07989__S _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__inv_2
X_11824_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11828_/C sky130_fd_sc_hd__nor2_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15592_/CLK _15592_/D _14661_/Y vssd1 vssd1 vccd1 vccd1 _15592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14543_/Y sky130_fd_sc_hd__inv_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11862_/B _11755_/B vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__xnor2_2
XFILLER_186_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08393__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10706_ _10706_/A _10706_/B _11012_/A vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__and3_1
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14474_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14474_/Y sky130_fd_sc_hd__inv_2
X_11686_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__or2_1
XFILLER_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _13425_/A _13425_/B _13425_/C vssd1 vssd1 vccd1 vccd1 _13426_/B sky130_fd_sc_hd__nand3_1
XFILLER_174_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10637_ _15269_/Q _15170_/Q vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12924__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _13356_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__xnor2_1
X_10568_ _10568_/A vssd1 vssd1 vccd1 vccd1 _15032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12307_ _12280_/A _12280_/B _12278_/A vssd1 vssd1 vccd1 vccd1 _12326_/A sky130_fd_sc_hd__o21a_2
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10499_ _15254_/Q _15287_/Q vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__or2_1
XFILLER_114_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13287_ _13287_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__or2_1
XFILLER_170_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15026_ _15221_/CLK _15026_/D _14063_/Y vssd1 vssd1 vccd1 vccd1 _15026_/Q sky130_fd_sc_hd__dfrtp_1
X_12238_ _12238_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12240_/C sky130_fd_sc_hd__xnor2_1
XFILLER_29_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12169_ _12110_/S _12178_/A _12042_/B vssd1 vssd1 vccd1 vccd1 _12169_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater781_A _15616_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 x_i_0[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14586__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__A1 _07720_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08400_ _08401_/A _08437_/A vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__xor2_1
X_09380_ _09380_/A vssd1 vssd1 vccd1 vccd1 _15144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08331_ _11435_/A _08330_/Y _08263_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08331_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _08292_/B vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__inv_2
XFILLER_36_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08193_ _08194_/A _08194_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12834__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08523__S _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A1 input241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput320 _15662_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[2] sky130_fd_sc_hd__buf_2
XFILLER_160_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput331 output331/A vssd1 vssd1 vccd1 vccd1 y_i_4[12] sky130_fd_sc_hd__buf_2
Xoutput342 output342/A vssd1 vssd1 vccd1 vccd1 y_i_4[7] sky130_fd_sc_hd__buf_2
Xoutput353 _15677_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[1] sky130_fd_sc_hd__buf_2
Xoutput364 output364/A vssd1 vssd1 vccd1 vccd1 y_i_6[11] sky130_fd_sc_hd__buf_2
Xoutput375 output375/A vssd1 vssd1 vccd1 vccd1 y_i_6[6] sky130_fd_sc_hd__buf_2
XFILLER_114_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput386 output386/A vssd1 vssd1 vccd1 vccd1 y_i_7[16] sky130_fd_sc_hd__buf_2
Xoutput397 output397/A vssd1 vssd1 vccd1 vccd1 y_r_0[10] sky130_fd_sc_hd__buf_2
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_578 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07977_ _15797_/Q vssd1 vssd1 vccd1 vccd1 _11678_/A sky130_fd_sc_hd__buf_6
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09716_ _09716_/A _09716_/B vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_751 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09647_ _09645_/A _09645_/B _09646_/X vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14496__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11913__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _15438_/Q _15422_/Q vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__nor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07602__S _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08529_ _08697_/B _08529_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11540_ _11828_/A _11827_/C _11828_/B vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__and3_1
XFILLER_195_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11471_ _12312_/S _11471_/B vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__nand2_1
XFILLER_183_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input195_A x_r_4[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12744__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13210_ _13210_/A _13715_/A vssd1 vssd1 vccd1 vccd1 _13563_/B sky130_fd_sc_hd__xor2_4
X_10422_ _10421_/A _10421_/C _10421_/B vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__a21oi_1
XFILLER_167_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14190_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10353_ _10352_/A _10352_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__a21o_1
X_13141_ _13712_/A _13712_/B _13713_/B _13703_/B _13133_/B vssd1 vssd1 vccd1 vccd1
+ _13210_/A sky130_fd_sc_hd__a32o_2
XFILLER_164_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ _13072_/A _13072_/B vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input56_A x_i_3[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _15084_/Q _15249_/Q vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__or2b_1
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12023_ _12099_/B _12023_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__and2_1
XFILLER_133_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10711__B _15282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13974_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13974_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15713_ _15791_/CLK _15713_/D _14789_/Y vssd1 vssd1 vccd1 vccd1 _15713_/Q sky130_fd_sc_hd__dfrtp_1
X_12925_ _13422_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07702__A1 _07702_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15644_ _15679_/CLK _15644_/D _14716_/Y vssd1 vssd1 vccd1 vccd1 _15644_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12856_ _12959_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12638__B _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07512__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _12055_/A _11523_/B _11977_/A vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15575_ _15575_/CLK _15575_/D _14644_/Y vssd1 vssd1 vccd1 vccd1 _15575_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12787_ _12787_/A _12787_/B vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__xnor2_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14526_/A vssd1 vssd1 vccd1 vccd1 _14526_/Y sky130_fd_sc_hd__inv_2
X_11738_ _11922_/B _11738_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__nor2_1
XFILLER_187_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1005 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14457_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14457_/Y sky130_fd_sc_hd__inv_2
X_11669_ _11898_/A vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__inv_2
XANTENNA__12654__A _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater627_A _11357_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ _13404_/Y _13574_/A _13407_/X vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__o21a_1
X_14388_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14388_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07769__A1 input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_712 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13339_ _13340_/A _13340_/B _13340_/C vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__a21o_1
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15009_ _15175_/CLK _15009_/D _14045_/Y vssd1 vssd1 vccd1 vccd1 _15009_/Q sky130_fd_sc_hd__dfrtp_1
X_07900_ _15317_/Q input131/X _07900_/S vssd1 vssd1 vccd1 vccd1 _07901_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08880_ _08950_/A _08877_/B _08879_/X vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07831_ _07831_/A vssd1 vssd1 vccd1 vccd1 _15352_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater801 _15590_/Q vssd1 vssd1 vccd1 vccd1 repeater801/X sky130_fd_sc_hd__buf_2
XFILLER_96_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater812 _15577_/Q vssd1 vssd1 vccd1 vccd1 repeater812/X sky130_fd_sc_hd__buf_2
XFILLER_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater823 input92/X vssd1 vssd1 vccd1 vccd1 _07471_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater834 input83/X vssd1 vssd1 vccd1 vccd1 _07477_/A1 sky130_fd_sc_hd__buf_4
XFILLER_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater845 input62/X vssd1 vssd1 vccd1 vccd1 repeater845/X sky130_fd_sc_hd__buf_2
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07762_ _07762_/A vssd1 vssd1 vccd1 vccd1 _15386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater856 input54/X vssd1 vssd1 vccd1 vccd1 _07420_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater867 input35/X vssd1 vssd1 vccd1 vccd1 _07575_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater878 input249/X vssd1 vssd1 vccd1 vccd1 _07642_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater889 input235/X vssd1 vssd1 vccd1 vccd1 repeater889/X sky130_fd_sc_hd__buf_2
X_09501_ _09501_/A _09501_/B vssd1 vssd1 vccd1 vccd1 _15254_/D sky130_fd_sc_hd__xnor2_1
X_07693_ _15419_/Q input191/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07694_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07930__B _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _15531_/Q _15515_/Q vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07422__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _15401_/Q _15385_/Q vssd1 vssd1 vccd1 vccd1 _09363_/X sky130_fd_sc_hd__and2b_1
XFILLER_52_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ _08324_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08314_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09294_ _15402_/Q _15386_/Q vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ _08265_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08279_/A sky130_fd_sc_hd__xnor2_2
XFILLER_193_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__xnor2_1
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15297__D _15297_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_63_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09873__A _15187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_121_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _15007_/D sky130_fd_sc_hd__xor2_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12739__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15760__D _15760_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _12710_/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input110_A x_i_6[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input208_A x_r_4[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ _13690_/A _13690_/B vssd1 vssd1 vccd1 vccd1 _13690_/X sky130_fd_sc_hd__or2_1
XFILLER_71_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_136_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ _15051_/Q _12711_/B vssd1 vssd1 vccd1 vccd1 _12718_/B sky130_fd_sc_hd__xnor2_1
XFILLER_19_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15360_ _15722_/CLK _15360_/D _14415_/Y vssd1 vssd1 vccd1 vccd1 _15360_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12572_ _12340_/A _12571_/B _12340_/B vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__a21bo_1
XFILLER_157_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14311_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14311_/Y sky130_fd_sc_hd__inv_2
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__xor2_1
XFILLER_7_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15291_ _15553_/CLK _15291_/D _14343_/Y vssd1 vssd1 vccd1 vccd1 _15291_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14242_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14242_/Y sky130_fd_sc_hd__inv_2
X_11454_ _11531_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__xnor2_1
XFILLER_184_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _14945_/D sky130_fd_sc_hd__xor2_1
X_14173_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14173_/Y sky130_fd_sc_hd__inv_2
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__xor2_4
XFILLER_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07620__A0 _15455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _13124_/A _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__and3_1
X_10336_ _10467_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _15784_/D sky130_fd_sc_hd__xnor2_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _12973_/A _13051_/Y _13057_/C _13053_/X _13054_/Y vssd1 vssd1 vccd1 vccd1
+ _13058_/A sky130_fd_sc_hd__a221oi_2
X_10267_ _10267_/A _10267_/B _11418_/A vssd1 vssd1 vccd1 vccd1 _10267_/X sky130_fd_sc_hd__and3_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12006_ _12062_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12008_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10198_ _10197_/A _10197_/B _11394_/A vssd1 vssd1 vccd1 vccd1 _10199_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_output427_A output427/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13957_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13957_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_924 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11553__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12908_ _12909_/B _13018_/B _13020_/A vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__a21o_2
XFILLER_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _15059_/D sky130_fd_sc_hd__xor2_1
XFILLER_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15627_ _15761_/CLK _15627_/D _14698_/Y vssd1 vssd1 vccd1 vccd1 _15627_/Q sky130_fd_sc_hd__dfrtp_1
X_12839_ _13021_/B _12913_/B vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__xor2_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14864__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater744_A _15656_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07439__A0 _15544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _15558_/CLK _15558_/D _14625_/Y vssd1 vssd1 vccd1 vccd1 _15559_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_72_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11699__S _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14509_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater911_A input202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15489_ _15664_/CLK _15489_/D _14552_/Y vssd1 vssd1 vccd1 vccd1 _15489_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08030_ _11447_/C _08097_/B _11435_/A vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__mux2_1
XFILLER_200_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 x_i_1[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_2
Xinput41 x_i_2[15] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
Xinput52 x_i_3[10] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
Xinput63 x_i_3[6] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_892 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput74 x_i_4[1] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput85 x_i_5[11] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput96 x_i_5[7] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09981_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _14927_/D sky130_fd_sc_hd__xnor2_1
XFILLER_192_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__A _11728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _08931_/Y _15459_/Q _08927_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07925__B _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _15465_/Q _15449_/Q vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08102__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater620 _11041_/Y vssd1 vssd1 vccd1 vccd1 repeater620/X sky130_fd_sc_hd__buf_2
Xrepeater631 _10733_/Y vssd1 vssd1 vccd1 vccd1 output406/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ _15360_/Q _07814_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07815_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13943__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater642 _11250_/X vssd1 vssd1 vccd1 vccd1 output472/A sky130_fd_sc_hd__clkbuf_2
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater653 _07966_/X vssd1 vssd1 vccd1 vccd1 repeater653/X sky130_fd_sc_hd__buf_2
X_08794_ _15341_/Q _15325_/Q vssd1 vssd1 vccd1 vccd1 _08795_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08898__B_N _15455_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater664 _14750_/A vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__buf_4
Xrepeater675 _14642_/X vssd1 vssd1 vccd1 vccd1 _14656_/A sky130_fd_sc_hd__clkbuf_8
X_07745_ _07745_/A vssd1 vssd1 vccd1 vccd1 _15394_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater686 _14376_/A vssd1 vssd1 vccd1 vccd1 _14369_/A sky130_fd_sc_hd__buf_6
Xrepeater697 _08290_/B vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__buf_6
XANTENNA__15580__D _15580_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07676_ _07676_/A vssd1 vssd1 vccd1 vccd1 _15428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _09414_/A _09414_/B _09498_/A vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14774__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09346_ _15411_/Q _15395_/Q _09345_/X vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__a21oi_2
XFILLER_205_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11910__B _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _15397_/Q _15381_/Q _09351_/C vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__a21oi_1
XFILLER_193_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ _08239_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08159_ _11687_/A vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__clkinv_2
XFILLER_134_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _15747_/Q _15025_/Q vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__or2_1
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _15140_/Q _15305_/Q vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14014__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input158_A x_r_1[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _15210_/Q _15111_/Q vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__nand2_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14860_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _13809_/A _13809_/B _13810_/X vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__o21a_2
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14791_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14791_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input19_A x_i_1[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07669__A0 _15431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ _14980_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__xor2_4
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10954_ _14968_/Q _10953_/Y _10952_/B vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__a21oi_4
XFILLER_95_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__B _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13673_ _14974_/Q _13820_/B vssd1 vssd1 vccd1 vccd1 _13819_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__14684__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _14959_/Q _14893_/Q vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15412_ _15575_/CLK _15412_/D _14471_/Y vssd1 vssd1 vccd1 vccd1 _15412_/Q sky130_fd_sc_hd__dfrtp_1
X_12624_ _15759_/Q vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__inv_2
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15343_ _15758_/CLK _15343_/D _14397_/Y vssd1 vssd1 vccd1 vccd1 _15343_/Q sky130_fd_sc_hd__dfrtp_1
X_12555_ _12556_/A _12556_/C _12556_/B vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__a21oi_1
XFILLER_157_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11506_ _12360_/B _11507_/B vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__or2_1
XFILLER_106_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15274_ _15279_/CLK _15274_/D _14325_/Y vssd1 vssd1 vccd1 vccd1 _15274_/Q sky130_fd_sc_hd__dfrtp_1
X_12486_ _12497_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__xnor2_2
XFILLER_184_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output377_A output377/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14225_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11437_ _08014_/A _08014_/B _11436_/X vssd1 vssd1 vccd1 vccd1 _11531_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08397__A1 _08396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14156_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11368_ _11191_/Y _11367_/B _11193_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__o21ai_4
XFILLER_4_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13107_ _13491_/S _13390_/A _13106_/C vssd1 vssd1 vccd1 vccd1 _13108_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10319_ _10317_/Y _10319_/B vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__and2b_2
XFILLER_140_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11299_ _11298_/A _11298_/B _10801_/B vssd1 vssd1 vccd1 vccd1 _11300_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13037_/Y _12959_/A _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _13040_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_504 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater694_A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14859__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater861_A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14989_ _15119_/CLK _14989_/D _14023_/Y vssd1 vssd1 vccd1 vccd1 _14989_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater959_A input136/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07530_ _15499_/Q input111/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07461_ _15533_/Q _07461_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14594__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _09200_/A _09667_/B vssd1 vssd1 vccd1 vccd1 _15296_/D sky130_fd_sc_hd__xor2_1
XFILLER_210_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07392_ _15571_/Q _07392_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07393_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07700__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ _09129_/A _09265_/A _09130_/Y vssd1 vssd1 vccd1 vccd1 _09133_/A sky130_fd_sc_hd__o21ai_1
XFILLER_175_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07832__A0 _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ _15379_/Q vssd1 vssd1 vccd1 vccd1 _09062_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08013_ _11436_/B _08013_/B vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_163_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13938__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11458__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _15233_/Q _15200_/Q vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__or2b_1
XFILLER_89_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08915_ _08914_/A _08914_/B _08967_/A vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09895_ _15222_/Q _15189_/Q vssd1 vssd1 vccd1 vccd1 _09896_/C sky130_fd_sc_hd__and2b_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14769__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _13914_/A _08844_/B _08845_/X vssd1 vssd1 vccd1 vccd1 _15085_/D sky130_fd_sc_hd__a21o_1
XFILLER_58_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _13880_/A _08772_/B _08776_/X vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14919__D _14919_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _15402_/Q input222/X _07750_/S vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__mux2_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07659_ _15436_/Q _07659_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _15276_/Q _15177_/Q vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__or2_1
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07610__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _15408_/Q _15392_/Q vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__and2_1
XFILLER_16_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14009__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12340_ _12340_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12571_/A sky130_fd_sc_hd__nand2_2
XFILLER_167_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _12271_/A vssd1 vssd1 vccd1 vccd1 _15589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14010_/Y sky130_fd_sc_hd__inv_2
X_11222_ _11222_/A _11230_/A vssd1 vssd1 vccd1 vccd1 _11379_/A sky130_fd_sc_hd__nand2_2
XFILLER_175_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13567__B _13567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11153_ _11153_/A _11153_/B _11355_/A vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__and3_1
XFILLER_161_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _15119_/Q vssd1 vssd1 vccd1 vccd1 _10104_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11084_ _11084_/A _11084_/B vssd1 vssd1 vccd1 vccd1 _11346_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11087__B _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput220 x_r_5[3] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14679__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput231 x_r_6[13] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__clkbuf_2
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _10395_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _14975_/D sky130_fd_sc_hd__xnor2_1
Xinput242 x_r_6[9] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14912_ _15532_/CLK _14912_/D _13942_/Y vssd1 vssd1 vccd1 vccd1 _14912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput253 x_r_7[4] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14843_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14843_/Y sky130_fd_sc_hd__inv_2
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08396__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14774_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _11986_/A _11986_/B vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__nand2_1
XFILLER_189_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11989__A2 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ _13725_/A _13725_/B _13725_/C vssd1 vssd1 vccd1 vccd1 _13841_/B sky130_fd_sc_hd__and3_1
XFILLER_56_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_866 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _10937_/A _10945_/A vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_899 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13656_ _13669_/A _13646_/B _13646_/C vssd1 vssd1 vccd1 vccd1 _13656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_143_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ _10867_/A _10867_/B _11107_/A vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output494_A output494/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12938__A1 _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _12607_/A _12607_/B vssd1 vssd1 vccd1 vccd1 _15688_/D sky130_fd_sc_hd__xor2_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _15773_/Q _13588_/B vssd1 vssd1 vccd1 vccd1 _13587_/Y sky130_fd_sc_hd__nand2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _15724_/Q _15790_/Q vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__and2b_1
XFILLER_200_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15326_ _15341_/CLK _15326_/D _14379_/Y vssd1 vssd1 vccd1 vccd1 _15326_/Q sky130_fd_sc_hd__dfrtp_1
X_12538_ _11725_/B _15730_/Q vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15257_ _15542_/CLK _15257_/D _14307_/Y vssd1 vssd1 vccd1 vccd1 _15257_/Q sky130_fd_sc_hd__dfrtp_1
X_12469_ _12484_/B _12475_/C _14949_/Q vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12662__A _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater707_A _07575_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14208_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15188_ _15192_/CLK _15188_/D _14233_/Y vssd1 vssd1 vccd1 vccd1 _15188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14139_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14158_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14589__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _13634_/B sky130_fd_sc_hd__xor2_4
X_09680_ _09680_/A _09680_/B vssd1 vssd1 vccd1 vccd1 _15315_/D sky130_fd_sc_hd__xnor2_1
XFILLER_95_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08631_ _08631_/A _08631_/B vssd1 vssd1 vccd1 vccd1 _08631_/X sky130_fd_sc_hd__and2_1
XFILLER_82_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08562_ _08598_/A _08597_/A vssd1 vssd1 vccd1 vccd1 _08566_/C sky130_fd_sc_hd__or2_1
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ _07513_/A vssd1 vssd1 vccd1 vccd1 _15508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ _12871_/A _12780_/A vssd1 vssd1 vccd1 vccd1 _08496_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07444_ _07444_/A vssd1 vssd1 vccd1 vccd1 _15542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07430__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09114_ _09114_/A _09250_/A _09114_/C vssd1 vssd1 vccd1 vccd1 _09116_/A sky130_fd_sc_hd__nor3_1
XANTENNA__11601__A1 _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_924 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09270__A2 _15491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09045_ _09045_/A _09045_/B _13622_/A vssd1 vssd1 vccd1 vccd1 _09045_/X sky130_fd_sc_hd__and3_1
XFILLER_190_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_92 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09947_ _09946_/A _09946_/B _09997_/A vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14499__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _15188_/Q _15221_/Q vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__or2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08497__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08829_ _15330_/Q _15346_/Q vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__and2b_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _12254_/A _12144_/A _11839_/C vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__a21oi_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10569__B_N _15297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11771_ _11876_/A _11667_/B _11672_/B _11770_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12747__A _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13510_ _13510_/A _13791_/B vssd1 vssd1 vccd1 vccd1 _13588_/B sky130_fd_sc_hd__xor2_2
XFILLER_53_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10722_ _10722_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _10723_/B sky130_fd_sc_hd__and2_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11840__A1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14490_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13441_ _13441_/A _13441_/B _13441_/C vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__and3_1
X_10653_ _10645_/Y _10649_/B _10647_/B vssd1 vssd1 vccd1 vccd1 _10654_/B sky130_fd_sc_hd__o21ai_4
XFILLER_142_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13593__A1 _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input86_A x_i_5[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _13372_/A _13372_/B vssd1 vssd1 vccd1 vccd1 _13399_/A sky130_fd_sc_hd__xor2_1
XFILLER_10_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10584_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10585_/B sky130_fd_sc_hd__and2_1
XFILLER_155_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15111_ _15375_/CLK _15111_/D _14152_/Y vssd1 vssd1 vccd1 vccd1 _15111_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _15740_/Q _12323_/B vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__and2_1
XFILLER_182_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _15467_/CLK _15042_/D _14080_/Y vssd1 vssd1 vccd1 vccd1 _15042_/Q sky130_fd_sc_hd__dfrtp_1
X_12254_ _12254_/A _12254_/B vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__xnor2_1
XFILLER_177_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ _15029_/Q _15751_/Q vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__or2b_1
X_12185_ _12185_/A _12185_/B vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__xnor2_2
XFILLER_150_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _11134_/A _11134_/B _11135_/X vssd1 vssd1 vccd1 vccd1 _11137_/B sky130_fd_sc_hd__a21o_2
XFILLER_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_683 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _11335_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/Y sky130_fd_sc_hd__xnor2_1
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14202__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11545__B _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _15203_/Q _15104_/Q vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__nand2_1
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output507_A output507/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14826_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12069__D1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14757_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14757_/Y sky130_fd_sc_hd__inv_2
X_11969_ _12046_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__or2_1
XFILLER_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_137_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15532_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08854__B _15447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _13708_/A _13830_/B vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__nor2_1
X_14688_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14688_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ _13639_/A _13639_/B vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_repeater824_A input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_740 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14872__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15309_ _15568_/CLK _15309_/D _14362_/Y vssd1 vssd1 vccd1 vccd1 _15309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10905__A _10905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput502 _11233_/X vssd1 vssd1 vccd1 vccd1 y_r_6[13] sky130_fd_sc_hd__buf_2
XFILLER_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput513 output513/A vssd1 vssd1 vccd1 vccd1 y_r_6[8] sky130_fd_sc_hd__buf_2
XFILLER_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput524 output524/A vssd1 vssd1 vccd1 vccd1 y_r_7[2] sky130_fd_sc_hd__buf_2
XFILLER_160_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13887__A2 _15322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13000__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09801_ _09801_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _15163_/D sky130_fd_sc_hd__nor2_1
XFILLER_99_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07993_ _15804_/Q vssd1 vssd1 vccd1 vccd1 _12178_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_68_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11736__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _15062_/Q _15095_/Q _09728_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10640__A _15270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_985 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09663_ _09663_/A _09663_/B _09663_/C vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__and3_1
XFILLER_41_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13951__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _08728_/A _12970_/A vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__or2_1
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09594_ _15424_/Q _15440_/Q vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__or2b_1
XFILLER_199_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08545_ _08558_/A _08566_/A _08566_/B vssd1 vssd1 vccd1 vccd1 _08551_/A sky130_fd_sc_hd__or3_1
XFILLER_23_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_128_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11471__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_392 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08476_ _08478_/B _08728_/A _08478_/A vssd1 vssd1 vccd1 vccd1 _08552_/A sky130_fd_sc_hd__or3b_1
XFILLER_210_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ _07427_/A vssd1 vssd1 vccd1 vccd1 _15550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ _15359_/Q _15375_/Q vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__or2b_1
XFILLER_156_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input140_A x_r_0[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13990_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14022__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input238_A x_r_6[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _12900_/A _12900_/B _12940_/Y vssd1 vssd1 vccd1 vccd1 _12943_/B sky130_fd_sc_hd__o21a_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15660_ _15663_/CLK _15660_/D _14733_/Y vssd1 vssd1 vccd1 vccd1 _15660_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12872_/A _12802_/A vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__or2b_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14611_/Y sky130_fd_sc_hd__inv_2
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11825_/B _11779_/B vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__or2b_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15648_/CLK _15591_/D _14660_/Y vssd1 vssd1 vccd1 vccd1 _15591_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_119_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15347_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14542_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11754_ _11714_/A _11714_/B _11710_/A vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10705_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__nor2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14473_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11685_ _11685_/A _11685_/B vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__14692__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ _13425_/A _13425_/B _13425_/C vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__a21o_1
XFILLER_179_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10636_ _15269_/Q _15170_/Q vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12924__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ _15051_/Q _13355_/B vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__xnor2_1
X_10567_ _10565_/X _10572_/B vssd1 vssd1 vccd1 vccd1 _10568_/A sky130_fd_sc_hd__and2b_1
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ _15740_/Q vssd1 vssd1 vccd1 vccd1 _12319_/A sky130_fd_sc_hd__inv_2
XFILLER_182_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _13565_/A _13286_/B vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__xnor2_1
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10498_ _10498_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _15022_/D sky130_fd_sc_hd__nor2_1
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output457_A _15597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15025_ _15221_/CLK _15025_/D _14062_/Y vssd1 vssd1 vccd1 vccd1 _15025_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12237_ _12237_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12238_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ _12236_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__or2_1
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_749 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11556__A _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__B _15462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _11119_/A _11119_/B vssd1 vssd1 vccd1 vccd1 _11119_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12099_ _12099_/A _12099_/B _12553_/A vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__and3_1
XFILLER_110_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 x_i_0[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater774_A _15624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14867__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14809_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14809_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater941_A input160/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15789_ _15791_/CLK _15789_/D _14869_/Y vssd1 vssd1 vccd1 vccd1 _15789_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08330_ _11467_/A vssd1 vssd1 vccd1 vccd1 _08330_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11804__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08261_ _08265_/C _08257_/A _08257_/B _08277_/A _08277_/B vssd1 vssd1 vccd1 vccd1
+ _08279_/B sky130_fd_sc_hd__a32o_1
XFILLER_177_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ _08192_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08194_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14107__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13011__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput310 _10918_/X vssd1 vssd1 vccd1 vccd1 y_i_2[9] sky130_fd_sc_hd__buf_2
XFILLER_10_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput321 output321/A vssd1 vssd1 vccd1 vccd1 y_i_3[3] sky130_fd_sc_hd__buf_2
XFILLER_195_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput332 _11346_/X vssd1 vssd1 vccd1 vccd1 y_i_4[13] sky130_fd_sc_hd__buf_2
XFILLER_126_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13946__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A_N _15338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput343 output343/A vssd1 vssd1 vccd1 vccd1 y_i_4[8] sky130_fd_sc_hd__buf_2
XFILLER_161_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput354 output354/A vssd1 vssd1 vccd1 vccd1 y_i_5[2] sky130_fd_sc_hd__buf_2
Xoutput365 output365/A vssd1 vssd1 vccd1 vccd1 y_i_6[12] sky130_fd_sc_hd__buf_2
Xoutput376 _11117_/Y vssd1 vssd1 vccd1 vccd1 y_i_6[7] sky130_fd_sc_hd__buf_2
XFILLER_160_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput387 output387/A vssd1 vssd1 vccd1 vccd1 y_i_7[1] sky130_fd_sc_hd__buf_2
XFILLER_82_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput398 output398/A vssd1 vssd1 vccd1 vccd1 y_r_0[11] sky130_fd_sc_hd__buf_2
XFILLER_43_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15583__D _15583_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__B _15318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _15793_/Q vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__buf_4
X_09715_ _15060_/Q _15093_/Q vssd1 vssd1 vccd1 vccd1 _09716_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11185__B _15027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14777__A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _15567_/Q _15547_/Q vssd1 vssd1 vccd1 vccd1 _09646_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09577_ _09791_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _15176_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08529_/B sky130_fd_sc_hd__xnor2_1
XFILLER_208_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07475__A1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _08459_/A _08459_/B vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__xor2_1
XFILLER_169_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11470_ _11480_/A _11468_/Y _08162_/B _11469_/Y vssd1 vssd1 vccd1 vccd1 _11563_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12744__B _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ _10421_/A _10421_/B _10421_/C vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__and3_1
XFILLER_109_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input188_A x_r_3[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14017__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08975__A1 _15475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _15766_/Q vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__inv_2
X_10352_ _10352_/A _10352_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _10352_/X sky130_fd_sc_hd__and3_1
XFILLER_109_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08015__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _13071_/A vssd1 vssd1 vccd1 vccd1 _13072_/B sky130_fd_sc_hd__inv_2
X_10283_ _15083_/Q _10282_/Y _10281_/B vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08727__A1 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12022_ _12022_/A _12022_/B _12550_/A vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__nand3_1
XFILLER_183_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13575__B _13576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input49_A x_i_2[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13973_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13973_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14687__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15712_ _15712_/CLK _15712_/D _14788_/Y vssd1 vssd1 vccd1 vccd1 _15712_/Q sky130_fd_sc_hd__dfrtp_1
X_12924_ _13366_/A _13273_/A vssd1 vssd1 vccd1 vccd1 _12927_/A sky130_fd_sc_hd__nand2_1
XFILLER_47_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15643_ _15679_/CLK _15643_/D _14715_/Y vssd1 vssd1 vccd1 vccd1 _15643_/Q sky130_fd_sc_hd__dfrtp_2
X_12855_ _13381_/B _13220_/A _12854_/C vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__a21oi_1
XFILLER_62_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11898_/A _11876_/A _11806_/C vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__and3_1
XFILLER_15_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15574_ _15576_/CLK _15574_/D _14643_/Y vssd1 vssd1 vccd1 vccd1 _15574_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12787_/B sky130_fd_sc_hd__xnor2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14525_/Y sky130_fd_sc_hd__inv_2
X_11737_ _12204_/A _12088_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _11738_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14456_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14456_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11668_ _11898_/A _12055_/A _11668_/C vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__and3_1
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15668__D _15668_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ _13576_/B _15769_/Q vssd1 vssd1 vccd1 vccd1 _13407_/X sky130_fd_sc_hd__or2b_1
XFILLER_174_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10619_ _10619_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _15000_/D sky130_fd_sc_hd__xor2_1
X_14387_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14387_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11599_ _11599_/A _11668_/C vssd1 vssd1 vccd1 vccd1 _11600_/C sky130_fd_sc_hd__xnor2_1
XFILLER_31_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13338_ _13393_/B _13338_/B vssd1 vssd1 vccd1 vccd1 _13340_/C sky130_fd_sc_hd__nand2_1
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _13308_/B _13269_/B vssd1 vssd1 vccd1 vccd1 _13270_/C sky130_fd_sc_hd__or2_1
XFILLER_170_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15008_ _15008_/CLK _15008_/D _14044_/Y vssd1 vssd1 vccd1 vccd1 _15008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater891_A input233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11286__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07830_ _15352_/Q _07830_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07831_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater802 _15588_/Q vssd1 vssd1 vccd1 vccd1 output415/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater813 _15560_/Q vssd1 vssd1 vccd1 vccd1 output259/A sky130_fd_sc_hd__buf_4
XFILLER_116_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater824 input91/X vssd1 vssd1 vccd1 vccd1 _07473_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater835 input81/X vssd1 vssd1 vccd1 vccd1 _07591_/A1 sky130_fd_sc_hd__clkbuf_2
X_07761_ _15386_/Q _07761_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__mux2_1
Xrepeater846 repeater847/X vssd1 vssd1 vccd1 vccd1 _07437_/A1 sky130_fd_sc_hd__buf_4
Xrepeater857 input53/X vssd1 vssd1 vccd1 vccd1 _07422_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14597__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater868 repeater869/X vssd1 vssd1 vccd1 vccd1 _07494_/A1 sky130_fd_sc_hd__buf_4
X_09500_ _15527_/Q _15511_/Q _09499_/X vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__a21o_1
Xrepeater879 input248/X vssd1 vssd1 vccd1 vccd1 _07644_/A1 sky130_fd_sc_hd__clkbuf_2
X_07692_ _07692_/A vssd1 vssd1 vccd1 vccd1 _15420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _15531_/Q _15515_/Q vssd1 vssd1 vccd1 vccd1 _09431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ _09362_/A _09362_/B vssd1 vssd1 vccd1 vccd1 _15139_/D sky130_fd_sc_hd__xor2_1
XFILLER_162_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08313_ _08276_/Y _08277_/Y _08314_/B _08324_/A _08312_/X vssd1 vssd1 vccd1 vccd1
+ _08313_/Y sky130_fd_sc_hd__a221oi_2
XANTENNA__07457__A1 _07457_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _15402_/Q _15386_/Q vssd1 vssd1 vccd1 vccd1 _09293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08244_ _08265_/B _08265_/C vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__nand2_1
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12564__B _12564_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08175_ _08175_/A _08174_/X vssd1 vssd1 vccd1 vccd1 _08176_/B sky130_fd_sc_hd__or2b_1
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07959_ _15251_/Q vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__clkinv_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10970_ _15269_/Q _10969_/Y _10968_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__a21o_1
XFILLER_71_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14300__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _09631_/C _09629_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__and2_1
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12640_ _12640_/A _12813_/C vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input103_A x_i_6[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12571_ _12571_/A _12571_/B vssd1 vssd1 vccd1 vccd1 _15625_/D sky130_fd_sc_hd__xor2_1
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_50_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15434_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14310_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14310_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11898_/A _12055_/A vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__xnor2_2
XFILLER_157_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _15553_/CLK _15290_/D _14342_/Y vssd1 vssd1 vccd1 vccd1 _15290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14241_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14241_/Y sky130_fd_sc_hd__inv_2
X_11453_ _11532_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A1 _15466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10404_ _15207_/Q _10403_/Y _10402_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__inv_2
X_11384_ _11382_/A _11382_/B _11383_/X vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__a21o_2
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13123_ _13123_/A vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__inv_2
X_10335_ _10327_/Y _10331_/B _10329_/B vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__07620__A1 _07620_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13054_/A _13054_/B vssd1 vssd1 vccd1 vccd1 _13054_/Y sky130_fd_sc_hd__nor2_1
X_10266_ _10266_/A _10274_/A vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__nand2_2
XFILLER_78_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12005_ _11924_/A _11924_/B _11921_/A vssd1 vssd1 vccd1 vccd1 _12006_/B sky130_fd_sc_hd__o21ai_1
XFILLER_121_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10197_ _10197_/A _10197_/B _11394_/A vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__and3_1
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output322_A _15664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14210__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13956_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13956_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11553__B _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__A1 input194/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _12985_/C _12907_/B vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__nand2_1
X_13887_ _15338_/Q _15322_/Q _13886_/X vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ _15741_/CLK _15626_/D _14697_/Y vssd1 vssd1 vccd1 vccd1 _15626_/Q sky130_fd_sc_hd__dfrtp_1
X_12838_ _13022_/A _12733_/B _13022_/B _12730_/A vssd1 vssd1 vccd1 vccd1 _12913_/B
+ sky130_fd_sc_hd__a31o_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07439__A1 _07439_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15557_ _15558_/CLK input1/X _14624_/Y vssd1 vssd1 vccd1 vccd1 _15558_/D sky130_fd_sc_hd__dfrtp_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12769_/A _13645_/B vssd1 vssd1 vccd1 vccd1 _12771_/A sky130_fd_sc_hd__or2_1
XANTENNA_repeater737_A _15665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12665__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15795_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__B _15449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14508_/Y sky130_fd_sc_hd__inv_2
X_15488_ _15511_/CLK _15488_/D _14551_/Y vssd1 vssd1 vccd1 vccd1 _15488_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput20 x_i_1[10] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater904_A input215/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14439_/Y sky130_fd_sc_hd__inv_2
Xinput31 x_i_1[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_2
XANTENNA__14880__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput42 x_i_2[1] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 x_i_3[11] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput64 x_i_3[7] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput75 x_i_4[2] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
Xinput86 x_i_5[12] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput97 x_i_5[8] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_2
XFILLER_196_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09980_ _09894_/A _09979_/B _09894_/B vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__a21boi_1
XFILLER_143_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08931_ _15475_/Q vssd1 vssd1 vccd1 vccd1 _08931_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _15465_/Q _15449_/Q vssd1 vssd1 vccd1 vccd1 _08862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater610 _11115_/Y vssd1 vssd1 vccd1 vccd1 output375/A sky130_fd_sc_hd__clkbuf_2
Xrepeater621 _10883_/Y vssd1 vssd1 vccd1 vccd1 output305/A sky130_fd_sc_hd__clkbuf_2
X_07813_ _07813_/A vssd1 vssd1 vccd1 vccd1 _15361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater632 repeater633/X vssd1 vssd1 vccd1 vccd1 output439/A sky130_fd_sc_hd__buf_4
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _15341_/Q _15325_/Q vssd1 vssd1 vccd1 vccd1 _08793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater643 _11149_/X vssd1 vssd1 vccd1 vccd1 output506/A sky130_fd_sc_hd__clkbuf_2
Xrepeater654 _07957_/X vssd1 vssd1 vccd1 vccd1 output294/A sky130_fd_sc_hd__clkbuf_2
Xrepeater665 _14753_/A vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__buf_6
X_07744_ _15394_/Q _07744_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07745_/A sky130_fd_sc_hd__mux2_1
Xrepeater676 _14559_/A vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__buf_6
XFILLER_84_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater687 _14376_/A vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__buf_4
XFILLER_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater698 _07795_/S vssd1 vssd1 vccd1 vccd1 _07765_/S sky130_fd_sc_hd__buf_4
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07675_ _15428_/Q _07675_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09414_ _09414_/A _09414_/B _09498_/A vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__nor3_1
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09419__A2 _15511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _15411_/Q _15395_/Q _09340_/A vssd1 vssd1 vccd1 vccd1 _09345_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15394_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_205_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09276_ _09354_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _09351_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08227_ _08239_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08237_/A sky130_fd_sc_hd__xor2_1
XFILLER_193_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07850__A1 _07850_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14790__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08158_ _11832_/A _11687_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__and3_1
XFILLER_180_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14940__D _14940_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07602__A1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _08094_/A _08076_/C _11806_/C vssd1 vssd1 vccd1 vccd1 _08090_/B sky130_fd_sc_hd__o21ai_1
XFILLER_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ _15140_/Q _15305_/Q vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__or2_1
XFILLER_122_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07608__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_99_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15752_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ _15210_/Q _15111_/Q vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__or2_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input220_A x_r_5[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _13810_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13810_/X sky130_fd_sc_hd__or2_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14790_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14030__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__A1 _07669_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ _13741_/A _13741_/B vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__nor2_2
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09124__A _15505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _14902_/Q vssd1 vssd1 vccd1 vccd1 _10953_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13672_ _13672_/A _13672_/B vssd1 vssd1 vccd1 vccd1 _13820_/B sky130_fd_sc_hd__xor2_4
XFILLER_71_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10884_ _14959_/Q _14893_/Q vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__or2_1
XFILLER_16_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15411_ _15411_/CLK _15411_/D _14470_/Y vssd1 vssd1 vccd1 vccd1 _15411_/Q sky130_fd_sc_hd__dfrtp_4
X_12623_ _15726_/Q _12623_/B vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__or2_1
XFILLER_188_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15809_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ _15752_/CLK _15342_/D _14396_/Y vssd1 vssd1 vccd1 vccd1 _15342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ _12549_/A _12550_/A _12549_/B _12098_/A _12551_/X vssd1 vssd1 vccd1 vccd1
+ _12556_/C sky130_fd_sc_hd__a311o_1
XFILLER_12_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _11431_/A _11431_/B _12525_/B _11504_/Y vssd1 vssd1 vccd1 vccd1 _11580_/A
+ sky130_fd_sc_hd__o31ai_2
X_15273_ _15592_/CLK _15273_/D _14324_/Y vssd1 vssd1 vccd1 vccd1 _15273_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _12485_/A _12485_/B vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__or2_1
XFILLER_145_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14224_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14224_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11436_ _08013_/B _11436_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__and2b_1
XFILLER_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output272_A output272/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08397__A2 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14155_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14155_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_98_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14205__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _13491_/S _13390_/A _13106_/C vssd1 vssd1 vccd1 vccd1 _13235_/B sky130_fd_sc_hd__and3_1
XANTENNA__07518__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10318_ _15125_/Q _15158_/Q vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14086_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14086_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08203__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ _11298_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__xor2_1
XFILLER_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13145_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _13037_/Y sky130_fd_sc_hd__nand2_1
X_10249_ _15243_/Q _15078_/Q vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__or2b_1
XFILLER_191_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15681__D _15681_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater687_A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1048 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_666 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14988_ _15119_/CLK _14988_/D _14022_/Y vssd1 vssd1 vccd1 vccd1 _14988_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater854_A repeater855/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14875__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07460_ _07460_/A vssd1 vssd1 vccd1 vccd1 _15534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08873__A _15467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15705_/CLK _15609_/D _14679_/Y vssd1 vssd1 vccd1 vccd1 _15609_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07391_ _07391_/A vssd1 vssd1 vccd1 vccd1 _15572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15498_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ _15506_/Q _15490_/Q vssd1 vssd1 vccd1 vccd1 _09130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_77_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09061_ _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _13631_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07832__A1 input171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ _08010_/Y _08052_/B _11584_/A vssd1 vssd1 vccd1 vccd1 _08013_/B sky130_fd_sc_hd__mux2_1
XFILLER_162_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07596__A0 _15467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14115__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07428__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _15200_/Q _15233_/Q vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_135_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13954__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _08914_/A _08914_/B _08967_/A vssd1 vssd1 vccd1 vccd1 _08914_/X sky130_fd_sc_hd__and3_1
XFILLER_134_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09894_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _15348_/Q _15332_/Q vssd1 vssd1 vccd1 vccd1 _08845_/X sky130_fd_sc_hd__and2b_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15591__D _15591_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11474__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08776_ _15336_/Q _15320_/Q vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__and2b_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _07727_/A vssd1 vssd1 vccd1 vccd1 _15403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07658_ _07658_/A vssd1 vssd1 vccd1 vccd1 _15437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07520__A0 _15504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_07589_ _15470_/Q input82/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09328_ _09328_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _15130_/D sky130_fd_sc_hd__xor2_4
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09258_/A _09258_/C _09258_/B vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ _12268_/X _12270_/B vssd1 vssd1 vccd1 vccd1 _12271_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ _15032_/Q _15754_/Q vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__or2b_1
XANTENNA_input170_A x_r_2[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07587__A0 _15471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14025__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _11150_/Y _11152_/B vssd1 vssd1 vccd1 vccd1 _11355_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09119__A _15504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10103_ _15284_/Q _10103_/B vssd1 vssd1 vccd1 vccd1 _10103_/Y sky130_fd_sc_hd__nand2_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11083_ _15000_/Q _14934_/Q vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__and2b_1
Xinput210 x_r_4[9] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_1
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input31_A x_i_1[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput221 x_r_5[4] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__clkbuf_1
Xinput232 x_r_6[14] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_2
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10034_ _10026_/Y _10030_/B _10028_/B vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__o21ai_1
X_14911_ _15532_/CLK _14911_/D _13941_/Y vssd1 vssd1 vccd1 vccd1 _14911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 x_r_7[0] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput254 x_r_7[5] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__clkbuf_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14861_/A sky130_fd_sc_hd__buf_8
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11985_ _11985_/A vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__inv_2
X_14773_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14773_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14695__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10936_ _14900_/Q _14966_/Q vssd1 vssd1 vccd1 vccd1 _10945_/A sky130_fd_sc_hd__or2b_1
X_13724_ _13725_/A _13725_/B _13725_/C vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__a21oi_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07801__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10867_ _10867_/A _10867_/B _11107_/A vssd1 vssd1 vccd1 vccd1 _10869_/A sky130_fd_sc_hd__and3_1
XFILLER_32_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13655_ _14973_/Q vssd1 vssd1 vccd1 vccd1 _13816_/A sky130_fd_sc_hd__clkinv_2
XFILLER_176_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08067__A1 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ _12601_/A _12604_/A _12601_/B _12605_/X vssd1 vssd1 vccd1 vccd1 _12607_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A _13586_/B vssd1 vssd1 vccd1 vccd1 _15609_/D sky130_fd_sc_hd__xnor2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _15723_/Q _15789_/Q _10797_/B vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__a21oi_4
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output487_A output487/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _12537_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _15614_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__07814__A1 _07814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15325_ _15341_/CLK _15325_/D _14378_/Y vssd1 vssd1 vccd1 vccd1 _15325_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ _12468_/A _12468_/B _12468_/C vssd1 vssd1 vccd1 vccd1 _12475_/C sky130_fd_sc_hd__nand3_1
X_15256_ _15542_/CLK _15256_/D _14306_/Y vssd1 vssd1 vccd1 vccd1 _15256_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14207_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14207_/Y sky130_fd_sc_hd__inv_2
X_11419_ _15081_/Q _15246_/Q vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__and2_1
XANTENNA_repeater602_A _11365_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ _15202_/CLK _15187_/D _14232_/Y vssd1 vssd1 vccd1 vccd1 _15187_/Q sky130_fd_sc_hd__dfrtp_1
X_12399_ _12410_/A _12399_/B vssd1 vssd1 vccd1 vccd1 _12400_/A sky130_fd_sc_hd__and2b_1
XFILLER_158_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14138_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14138_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14069_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14069_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_3_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15572_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08868__A _15466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__B _13790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater971_A input119/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08630_ _08564_/Y _08629_/X _08575_/B vssd1 vssd1 vccd1 vccd1 _08631_/B sky130_fd_sc_hd__a21bo_1
XFILLER_66_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07750__A0 _15391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ _13046_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08597_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07512_ _15508_/Q _07512_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07513_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08492_ _14916_/Q vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__buf_4
XFILLER_165_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07443_ _15542_/Q _07443_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07444_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09113_ _09113_/A _09113_/B vssd1 vssd1 vccd1 vccd1 _09114_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13949__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_936 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07947__A _15251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _09044_/A _09052_/A vssd1 vssd1 vccd1 vccd1 _13622_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10591__A1_N _15252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07569__A0 _15480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09946_ _09946_/A _09946_/B _09997_/A vssd1 vssd1 vccd1 vccd1 _09946_/X sky130_fd_sc_hd__and3_1
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _14956_/D sky130_fd_sc_hd__nor2_1
XFILLER_112_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08828_ _08828_/A vssd1 vssd1 vccd1 vccd1 _15081_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08759_ _15334_/Q _15318_/Q vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__and2b_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10721_ _10722_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__nor2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A2 _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13440_ _13441_/A _13441_/B _13441_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10652_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__nand2_2
XFILLER_41_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13371_ _13317_/A _13318_/A _13317_/B _13315_/A _13315_/B vssd1 vssd1 vccd1 vccd1
+ _13372_/B sky130_fd_sc_hd__o32a_1
XANTENNA__13593__A2 _15349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10583_ _15299_/Q _15266_/Q vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__or2b_1
XFILLER_103_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12322_ _12322_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _12322_/X sky130_fd_sc_hd__or2_1
XFILLER_10_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15110_ _15110_/CLK _15110_/D _14151_/Y vssd1 vssd1 vccd1 vccd1 _15110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input79_A x_i_4[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_766 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ _15509_/CLK _15041_/D _14078_/Y vssd1 vssd1 vccd1 vccd1 _15041_/Q sky130_fd_sc_hd__dfrtp_1
X_12253_ _12253_/A _12253_/B vssd1 vssd1 vccd1 vccd1 _12254_/B sky130_fd_sc_hd__nor2_1
XFILLER_142_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11204_ _11369_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11098__B _14936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ _12127_/A _12128_/A _12127_/B _12183_/X vssd1 vssd1 vccd1 vccd1 _12185_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_162_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _14967_/Q _14901_/Q vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__and2_1
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__nand2_1
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10017_ _15203_/Q _15104_/Q vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11545__C _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14825_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output402_A _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11842__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14756_/Y sky130_fd_sc_hd__inv_2
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ _11968_/A _11968_/B vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__and2_1
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ _14977_/Q vssd1 vssd1 vccd1 vccd1 _13708_/A sky130_fd_sc_hd__inv_2
XFILLER_189_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater552_A _10947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ _11121_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__nand2_1
X_11899_ _11980_/B _11899_/B vssd1 vssd1 vccd1 vccd1 _11901_/C sky130_fd_sc_hd__or2_1
X_14687_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14687_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _13638_/A _13638_/B vssd1 vssd1 vccd1 vccd1 _13639_/B sky130_fd_sc_hd__or2_2
XFILLER_158_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ _13564_/A _13566_/X _13564_/B _13567_/X vssd1 vssd1 vccd1 vccd1 _13570_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_200_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15308_ _15568_/CLK _15308_/D _14361_/Y vssd1 vssd1 vccd1 vccd1 _15308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput503 _11237_/Y vssd1 vssd1 vccd1 vccd1 y_r_6[14] sky130_fd_sc_hd__buf_2
X_15239_ _15472_/CLK _15239_/D _14288_/Y vssd1 vssd1 vccd1 vccd1 _15239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput514 _11203_/X vssd1 vssd1 vccd1 vccd1 y_r_6[9] sky130_fd_sc_hd__buf_2
Xoutput525 output525/A vssd1 vssd1 vccd1 vccd1 y_r_7[3] sky130_fd_sc_hd__buf_2
XFILLER_172_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08212__A1 _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09800_ _09799_/B _09799_/C _09799_/A vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__o21a_1
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07992_ _07990_/A _08087_/B _07991_/X vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__a21bo_1
XFILLER_86_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07706__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11736__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _09731_/A _09852_/A vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _09662_/A vssd1 vssd1 vccd1 vccd1 _15310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08613_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__and2_1
X_09593_ _09593_/A vssd1 vssd1 vccd1 vccd1 _15178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11752__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _13145_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _08566_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07441__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ _12803_/A _12688_/A vssd1 vssd1 vccd1 vccd1 _08478_/A sky130_fd_sc_hd__xor2_2
XFILLER_211_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07426_ _15550_/Q input66/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08780__B _15321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13398__B _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11199__A _15751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ _15374_/Q _15358_/Q vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__or2b_1
XFILLER_85_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11927__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14303__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07616__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09929_ _15195_/Q _15228_/Q vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__or2b_1
XFILLER_172_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _12940_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12940_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_input133_A x_r_0[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__xnor2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12758__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11662__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14610_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__inv_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11904_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11829_/A sky130_fd_sc_hd__nand2_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15717_/CLK _15590_/D _14659_/Y vssd1 vssd1 vccd1 vccd1 _15590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A _15507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _11863_/B _11753_/B vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__xor2_2
XFILLER_148_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14541_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__buf_6
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _15182_/Q _15281_/Q vssd1 vssd1 vccd1 vccd1 _10705_/B sky130_fd_sc_hd__and2b_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11684_ _11828_/A _11827_/C _11828_/B _11615_/A _11683_/X vssd1 vssd1 vccd1 vccd1
+ _11685_/B sky130_fd_sc_hd__a41o_1
XFILLER_186_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14472_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14472_/Y sky130_fd_sc_hd__inv_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10635_ _15268_/Q _15169_/Q _10634_/B vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__a21oi_4
XFILLER_139_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13423_ _13470_/B _13423_/B vssd1 vssd1 vccd1 vccd1 _13425_/C sky130_fd_sc_hd__nand2_1
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13355_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10566_ _10565_/A _10565_/B _10616_/A vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__a21o_1
XFILLER_155_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _12566_/A _12301_/B _12304_/Y vssd1 vssd1 vccd1 vccd1 _12321_/A sky130_fd_sc_hd__a21o_1
XFILLER_170_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13285_ _13211_/A _13563_/B _13409_/A vssd1 vssd1 vccd1 vccd1 _13286_/B sky130_fd_sc_hd__o21ai_1
X_10497_ _10496_/A _10496_/B _10592_/A vssd1 vssd1 vccd1 vccd1 _10498_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ _12236_/A _12236_/B _12236_/C vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__nor3_1
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15024_ _15221_/CLK _15024_/D _14061_/Y vssd1 vssd1 vccd1 vccd1 _15024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output352_A output352/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11837__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12167_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__and2_1
XANTENNA__14213__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07526__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ _10900_/A _11117_/B _10900_/B vssd1 vssd1 vccd1 vccd1 _11119_/B sky130_fd_sc_hd__a21boi_4
XFILLER_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12098_ _12098_/A _12556_/A vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__nor2b_2
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _11049_/A _11049_/B vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__nand2_2
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 x_i_0[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater767_A _15631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12668__A _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__B _15448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14808_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14808_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13254__A1 _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15788_ _15791_/CLK _15788_/D _14868_/Y vssd1 vssd1 vccd1 vccd1 _15788_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14739_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11804__A2 _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14883__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater934_A repeater935/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _08265_/C _08260_/B vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__xnor2_1
XFILLER_162_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _08209_/A _08209_/B _08190_/Y vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__a21oi_1
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput300 output300/A vssd1 vssd1 vccd1 vccd1 y_i_2[15] sky130_fd_sc_hd__buf_2
XFILLER_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput311 output311/A vssd1 vssd1 vccd1 vccd1 y_i_3[0] sky130_fd_sc_hd__buf_2
XFILLER_10_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput322 _15664_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[4] sky130_fd_sc_hd__buf_2
XFILLER_105_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput333 _11348_/X vssd1 vssd1 vccd1 vccd1 y_i_4[14] sky130_fd_sc_hd__buf_2
XFILLER_195_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput344 output344/A vssd1 vssd1 vccd1 vccd1 y_i_4[9] sky130_fd_sc_hd__buf_2
XFILLER_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput355 output355/A vssd1 vssd1 vccd1 vccd1 y_i_5[3] sky130_fd_sc_hd__buf_2
XFILLER_126_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput366 output366/A vssd1 vssd1 vccd1 vccd1 y_i_6[13] sky130_fd_sc_hd__buf_2
XFILLER_0_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput377 output377/A vssd1 vssd1 vccd1 vccd1 y_i_6[8] sky130_fd_sc_hd__buf_2
XANTENNA__10651__A _15272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput388 _15694_/Q vssd1 vssd1 vccd1 vccd1 y_i_7[2] sky130_fd_sc_hd__buf_2
XFILLER_114_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput399 _10782_/X vssd1 vssd1 vccd1 vccd1 y_r_0[12] sky130_fd_sc_hd__buf_2
XANTENNA__14123__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07975_ _07975_/A vssd1 vssd1 vccd1 vccd1 _07975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09714_ _15060_/Q _15093_/Q vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__or2_1
XANTENNA__13962__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09645_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _15306_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09788_/A _09571_/B _09575_/X vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__a21o_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__C _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12297__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10297__A2_N _15153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08528_/B sky130_fd_sc_hd__xor2_1
XFILLER_150_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14793__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _08458_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08459_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07409_ _07409_/A vssd1 vssd1 vccd1 vccd1 _15563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_839 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08389_ _08412_/A _08412_/B vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__xnor2_1
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10420_ _10420_/A vssd1 vssd1 vccd1 vccd1 _14948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08424__A1 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _10351_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__nor2_1
XFILLER_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13070_ _13070_/A vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__inv_2
XFILLER_152_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ _15248_/Q vssd1 vssd1 vccd1 vccd1 _10282_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12021_ _12022_/A _12022_/B _12550_/A vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08727__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input250_A x_r_7[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08031__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13972_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _15727_/CLK _15711_/D _14787_/Y vssd1 vssd1 vccd1 vccd1 _15711_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _12930_/B _12923_/B _12923_/C vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__or3_1
XFILLER_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ _15705_/CLK _15642_/D _14714_/Y vssd1 vssd1 vccd1 vccd1 _15642_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12039__A2 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ _13381_/B _13220_/A _12854_/C vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__and3_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_910 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11971_/B _11805_/B vssd1 vssd1 vccd1 vccd1 _11878_/A sky130_fd_sc_hd__nor2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15573_/CLK _15573_/D _14640_/Y vssd1 vssd1 vccd1 vccd1 _15573_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _08570_/A _12851_/B _12970_/A vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__mux2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14524_/Y sky130_fd_sc_hd__inv_2
X_11736_ _12204_/A _12088_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _11922_/B sky130_fd_sc_hd__and3_1
XFILLER_109_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14455_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14455_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11667_ _11876_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14208__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _13574_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _15637_/D sky130_fd_sc_hd__xnor2_4
X_10618_ _10616_/A _10616_/B _10617_/X vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08206__A _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _12122_/A _11977_/A vssd1 vssd1 vccd1 vccd1 _11668_/C sky130_fd_sc_hd__xor2_2
X_14386_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14386_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_850 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08966__A2 _15456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ _13381_/B _13337_/B vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__or2_1
X_10549_ _15294_/Q _15261_/Q vssd1 vssd1 vccd1 vccd1 _10558_/A sky130_fd_sc_hd__or2b_1
XFILLER_192_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268_ _13268_/A _13268_/B vssd1 vssd1 vccd1 vccd1 _13269_/B sky130_fd_sc_hd__nor2_1
XANTENNA__15684__D _15684_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11567__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _15008_/CLK _15007_/D _14043_/Y vssd1 vssd1 vccd1 vccd1 _15007_/Q sky130_fd_sc_hd__dfrtp_1
X_12219_ _12219_/A _12219_/B vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__xnor2_2
XFILLER_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _13197_/X _13274_/A vssd1 vssd1 vccd1 vccd1 _13201_/B sky130_fd_sc_hd__and2b_1
XFILLER_155_1062 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater803 _15587_/Q vssd1 vssd1 vccd1 vccd1 output414/A sky130_fd_sc_hd__buf_4
XANTENNA__14878__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater814 _15473_/Q vssd1 vssd1 vccd1 vccd1 _08968_/A sky130_fd_sc_hd__buf_2
Xrepeater825 input9/X vssd1 vssd1 vccd1 vccd1 _07610_/A1 sky130_fd_sc_hd__clkbuf_2
X_07760_ _07760_/A vssd1 vssd1 vccd1 vccd1 _15387_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clk/A sky130_fd_sc_hd__clkbuf_8
Xrepeater836 input77/X vssd1 vssd1 vccd1 vccd1 _07600_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater847 input61/X vssd1 vssd1 vccd1 vccd1 repeater847/X sky130_fd_sc_hd__buf_2
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater858 input47/X vssd1 vssd1 vccd1 vccd1 _07563_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11207__B_N _15752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater869 input33/X vssd1 vssd1 vccd1 vccd1 repeater869/X sky130_fd_sc_hd__buf_2
X_07691_ _15420_/Q input192/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ _09506_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _15272_/D sky130_fd_sc_hd__xor2_1
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09361_ _09359_/A _09359_/B _09360_/X vssd1 vssd1 vccd1 vccd1 _09362_/B sky130_fd_sc_hd__a21o_1
X_08312_ _08276_/Y _08277_/Y _08280_/Y _08342_/A _08311_/X vssd1 vssd1 vccd1 vccd1
+ _08312_/X sky130_fd_sc_hd__o221a_1
XFILLER_33_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ _09362_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _15123_/D sky130_fd_sc_hd__xnor2_1
XFILLER_61_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08243_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08265_/C sky130_fd_sc_hd__xor2_2
XFILLER_193_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10646__A _15271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__B _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14118__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ _08174_/A _08174_/B _08174_/C vssd1 vssd1 vccd1 vccd1 _08174_/X sky130_fd_sc_hd__or3_1
XFILLER_174_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13957__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14788__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07958_ _15152_/Q vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__inv_2
XFILLER_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13466__B2 _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ _07889_/A vssd1 vssd1 vccd1 vccd1 _15323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09628_ _15561_/Q _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__nand3_1
XFILLER_15_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _15433_/Q _15417_/Q vssd1 vssd1 vccd1 vccd1 _09559_/X sky130_fd_sc_hd__and2b_1
XFILLER_62_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12322_/X _12569_/B _12322_/A vssd1 vssd1 vccd1 vccd1 _12571_/B sky130_fd_sc_hd__o21ba_1
XFILLER_200_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ _11876_/A _11977_/A vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__A _15295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14028__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ _08023_/A _08023_/B _11451_/Y vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__a21oi_1
XFILLER_156_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14240_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14259_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_7_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ _15108_/Q vssd1 vssd1 vccd1 vccd1 _10403_/Y sky130_fd_sc_hd__inv_2
X_14171_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14171_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08948__A2 _15450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09070__A1 _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ _15755_/Q _15033_/Q vssd1 vssd1 vccd1 vccd1 _11383_/X sky130_fd_sc_hd__and2_1
XFILLER_178_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A x_i_3[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10341_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13122_ _13124_/A _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__a21o_1
XFILLER_180_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _12807_/Y _12804_/Y _13056_/B vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__o21a_1
X_10265_ _15246_/Q _15081_/Q vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__or2b_1
X_12004_ _12064_/A _12064_/B vssd1 vssd1 vccd1 vccd1 _12062_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10196_ _10194_/Y _10196_/B vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07384__A1 input120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14698__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08696__A _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13955_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13955_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output315_A _15673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12906_ _12906_/A _12906_/B _12906_/C vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__nand3_1
XFILLER_62_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _15338_/Q _15322_/Q _13885_/B vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15625_ _15717_/CLK _15625_/D _14696_/Y vssd1 vssd1 vccd1 vccd1 _15625_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12837_ _12835_/Y _12837_/B vssd1 vssd1 vccd1 vccd1 _13021_/B sky130_fd_sc_hd__nand2b_2
XFILLER_146_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08776__A_N _15336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15556_ _15575_/CLK _15556_/D _14623_/Y vssd1 vssd1 vccd1 vccd1 _15556_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12768_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__xnor2_1
XFILLER_188_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12665__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14507_/Y sky130_fd_sc_hd__inv_2
X_11719_ _12378_/B _11719_/B vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__and2_1
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater632_A repeater633/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15487_ _15506_/CLK _15487_/D _14550_/Y vssd1 vssd1 vccd1 vccd1 _15487_/Q sky130_fd_sc_hd__dfrtp_1
X_12699_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12699_/Y sky130_fd_sc_hd__inv_2
X_14438_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14438_/Y sky130_fd_sc_hd__inv_2
Xinput10 x_i_0[1] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 x_i_1[11] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 x_i_1[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 x_i_2[2] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12196__A1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 x_i_3[12] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput65 x_i_3[8] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14369_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput76 x_i_4[3] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput87 x_i_5[13] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
Xinput98 x_i_5[9] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ _08930_/A _08930_/B vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__nand2_1
XFILLER_170_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _08942_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _15204_/D sky130_fd_sc_hd__xor2_1
Xrepeater600 _10758_/Y vssd1 vssd1 vccd1 vccd1 output411/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07812_ _15361_/Q input166/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07813_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater611 repeater612/X vssd1 vssd1 vccd1 vccd1 output273/A sky130_fd_sc_hd__buf_4
X_08792_ _13890_/A _08792_/B vssd1 vssd1 vccd1 vccd1 _15076_/D sky130_fd_sc_hd__xor2_1
Xrepeater622 _10743_/Y vssd1 vssd1 vccd1 vccd1 output408/A sky130_fd_sc_hd__buf_4
Xrepeater633 _11355_/Y vssd1 vssd1 vccd1 vccd1 repeater633/X sky130_fd_sc_hd__buf_2
XANTENNA__14401__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater644 _10863_/X vssd1 vssd1 vccd1 vccd1 output302/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07714__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater655 _07957_/X vssd1 vssd1 vccd1 vccd1 _15812_/A sky130_fd_sc_hd__clkbuf_2
X_07743_ _07743_/A vssd1 vssd1 vccd1 vccd1 _15395_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater666 _14740_/A vssd1 vssd1 vccd1 vccd1 _14739_/A sky130_fd_sc_hd__buf_6
Xrepeater677 _14559_/A vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_38_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater688 _14269_/A vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__buf_8
XFILLER_26_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater699 _07803_/S vssd1 vssd1 vccd1 vccd1 _07791_/S sky130_fd_sc_hd__buf_6
X_07674_ _07674_/A vssd1 vssd1 vccd1 vccd1 _15429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09413_ _15527_/Q _15511_/Q vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__xnor2_1
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11760__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _09344_/A vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _09275_/A _15398_/Q vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__or2b_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ _12088_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08157_/A _11491_/A _11467_/A vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__and3_1
XFILLER_193_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12591__A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08088_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08101_/A sky130_fd_sc_hd__xor2_1
XFILLER_106_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_886 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _10408_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _14978_/D sky130_fd_sc_hd__xnor2_2
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14311__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07624__S _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A2 _15485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13740_ _13740_/A _13740_/B _13740_/C vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__and3_1
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10952_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input213_A x_r_5[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13671_ _13648_/A _13648_/B _13652_/B _13669_/Y _13670_/Y vssd1 vssd1 vccd1 vccd1
+ _13672_/B sky130_fd_sc_hd__a41o_2
X_10883_ _10883_/A _10883_/B vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__nor2_2
XFILLER_73_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15410_ _15411_/CLK _15410_/D _14469_/Y vssd1 vssd1 vccd1 vccd1 _15410_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _12622_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _15692_/D sky130_fd_sc_hd__xnor2_1
XFILLER_189_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_750 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ _15341_/CLK _15341_/D _14395_/Y vssd1 vssd1 vccd1 vccd1 _15341_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ _12553_/A _12553_/B vssd1 vssd1 vccd1 vccd1 _15619_/D sky130_fd_sc_hd__xor2_1
XFILLER_196_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11504_ _15727_/Q _12527_/B vssd1 vssd1 vccd1 vccd1 _11504_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15272_ _15399_/CLK _15272_/D _14323_/Y vssd1 vssd1 vccd1 vccd1 _15272_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12484_ _12484_/A _12484_/B _12484_/C vssd1 vssd1 vccd1 vccd1 _12485_/B sky130_fd_sc_hd__and3_1
XFILLER_185_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14223_/Y sky130_fd_sc_hd__inv_2
X_11435_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14154_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14154_/Y sky130_fd_sc_hd__inv_2
X_11366_ _11186_/A _11365_/B _11186_/B vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__a21boi_4
XFILLER_153_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output265_A _11095_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10317_ _15125_/Q _15158_/Q vssd1 vssd1 vccd1 vccd1 _10317_/Y sky130_fd_sc_hd__nor2_1
X_13105_ _13150_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13106_/C sky130_fd_sc_hd__and2_1
X_11297_ _11296_/A _11296_/B _10794_/B vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__a21o_1
X_14085_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14085_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13036_/A _13036_/B vssd1 vssd1 vccd1 vccd1 _13040_/A sky130_fd_sc_hd__xnor2_1
X_10248_ _11408_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__nand2_1
XANTENNA_output432_A output432/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10179_ _15149_/Q _15314_/Q _10178_/B vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__14221__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07534__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14987_ _15809_/CLK _14987_/D _14021_/Y vssd1 vssd1 vccd1 vccd1 _14987_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater582_A _11277_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13938_ _14889_/A vssd1 vssd1 vccd1 vccd1 _13957_/A sky130_fd_sc_hd__buf_12
XFILLER_19_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13869_ _13869_/A _13869_/B vssd1 vssd1 vccd1 vccd1 _15675_/D sky130_fd_sc_hd__xnor2_1
XFILLER_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater847_A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08873__B _15451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ _15705_/CLK _15608_/D _14678_/Y vssd1 vssd1 vccd1 vccd1 _15608_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_210_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ _15572_/Q _07390_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07391_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15539_ _15539_/CLK _15539_/D _14605_/Y vssd1 vssd1 vccd1 vccd1 _15539_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _15380_/Q _15364_/Q vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__or2_1
XFILLER_176_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08011_ _11658_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _08052_/B sky130_fd_sc_hd__xor2_1
XFILLER_190_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07596__A1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09962_ _15199_/Q _09961_/Y _09960_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__a21oi_2
XFILLER_131_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08913_ _08913_/A _08921_/A vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09893_ _15190_/Q _15223_/Q vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08844_ _13914_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _15084_/D sky130_fd_sc_hd__xnor2_1
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14131__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09225__A _15495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11474__B _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08775_ _08773_/Y _08775_/B vssd1 vssd1 vccd1 vccd1 _13883_/A sky130_fd_sc_hd__nand2b_1
XFILLER_27_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13970__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ _15403_/Q _07726_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__mux2_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07657_ _15437_/Q input257/X _07687_/S vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07520__A1 input101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__B _15323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07588_ _07588_/A vssd1 vssd1 vccd1 vccd1 _15471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_750 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _09327_/A _09390_/A vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__nand2_2
XFILLER_142_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09258_ _09258_/A _09258_/B _09258_/C vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__and3_1
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__xnor2_1
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14951__D _14951_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09189_ _09189_/A _09659_/A _09189_/C vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__nor3_1
XFILLER_193_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14306__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11220_ _15754_/Q _15032_/Q vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__or2b_1
XFILLER_175_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07587__A1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _15744_/Q _15022_/Q vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1057 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input163_A x_r_2[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ _10102_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _15793_/D sky130_fd_sc_hd__xnor2_2
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _14934_/Q _15000_/Q vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput200 x_r_4[14] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_2
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15782__D _15782_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 x_r_5[0] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput222 x_r_5[5] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__clkbuf_2
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _10033_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _15532_/CLK _14910_/D _13940_/Y vssd1 vssd1 vccd1 vccd1 _14910_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput233 x_r_6[15] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14041__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 x_r_7[10] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__clkbuf_2
Xinput255 x_r_7[6] vssd1 vssd1 vccd1 vccd1 input255/X sky130_fd_sc_hd__clkbuf_1
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A x_i_1[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _14841_/A vssd1 vssd1 vccd1 vccd1 _14841_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14772_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ _11926_/B _11984_/B vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__and2b_1
XFILLER_1_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13723_ _13723_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13725_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__09500__A2 _15511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ _14966_/Q _14900_/Q vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__or2b_1
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _13654_/A _13812_/A vssd1 vssd1 vccd1 vccd1 _15694_/D sky130_fd_sc_hd__xnor2_4
X_10866_ _10864_/Y _10866_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__and2b_2
XFILLER_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12605_ _12471_/B _12602_/X _12471_/A vssd1 vssd1 vccd1 vccd1 _12605_/X sky130_fd_sc_hd__a21bo_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13585_ _13585_/A _13585_/B vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__nand2_1
XFILLER_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _10797_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15768_/CLK _15324_/D _14377_/Y vssd1 vssd1 vccd1 vccd1 _15324_/Q sky130_fd_sc_hd__dfrtp_2
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output382_A output382/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15255_ _15527_/CLK _15255_/D _14305_/Y vssd1 vssd1 vccd1 vccd1 _15255_/Q sky130_fd_sc_hd__dfrtp_1
X_12467_ _12468_/B _12468_/C _12468_/A vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14216__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14206_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14206_/Y sky130_fd_sc_hd__inv_2
X_11418_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _15738_/D sky130_fd_sc_hd__xor2_2
X_15186_ _15202_/CLK _15186_/D _14231_/Y vssd1 vssd1 vccd1 vccd1 _15186_/Q sky130_fd_sc_hd__dfrtp_1
X_12398_ _12398_/A _12398_/B _12588_/A vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__or3_1
XFILLER_153_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14137_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14137_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11349_ _11348_/A _11348_/B _11092_/B vssd1 vssd1 vccd1 vccd1 _11350_/B sky130_fd_sc_hd__a21o_1
XFILLER_141_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14068_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater797_A _15594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__B _15450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _12985_/C _13016_/X _13017_/X _13018_/X vssd1 vssd1 vccd1 vccd1 _13023_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater964_A input128/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14886__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A1 _07750_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08560_ _08566_/B _08560_/B vssd1 vssd1 vccd1 vccd1 _08598_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07511_ _07511_/A vssd1 vssd1 vccd1 vccd1 _15509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08491_ _13381_/B _08491_/B vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07502__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07442_ _07442_/A vssd1 vssd1 vccd1 vccd1 _15543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09112_/A _09254_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12853__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09043_ _15377_/Q _15361_/Q vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__or2b_1
XFILLER_135_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_948 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14126__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13030__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07439__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07569__A1 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13965__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _09945_/A _09953_/A vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09875_/A _09875_/B _09973_/A vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__a21oi_1
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08825_/X _08832_/B vssd1 vssd1 vccd1 vccd1 _08828_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14796__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _15317_/Q vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__inv_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07709_ _07709_/A vssd1 vssd1 vccd1 vccd1 _15412_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14946__D _14946_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08689_/A _08689_/B vssd1 vssd1 vccd1 vccd1 _08689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10720_ _11251_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _11248_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10651_ _15272_/Q _15173_/Q vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _13370_/A _13370_/B vssd1 vssd1 vccd1 vccd1 _13372_/A sky130_fd_sc_hd__or2_1
X_10582_ _15266_/Q _15299_/Q vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__or2b_1
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15777__D _15777_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ _12321_/A _12569_/A vssd1 vssd1 vccd1 vccd1 _15591_/D sky130_fd_sc_hd__xnor2_2
XFILLER_177_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14036__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _15509_/CLK _15040_/D _14077_/Y vssd1 vssd1 vccd1 vccd1 _15040_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12252_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__nor3_1
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _11369_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11203_/X sky130_fd_sc_hd__xor2_4
X_12183_ _12183_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ _11134_/A _11134_/B vssd1 vssd1 vccd1 vccd1 _11134_/X sky130_fd_sc_hd__xor2_4
XFILLER_27_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ _14930_/Q _14996_/Q _11061_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__a21o_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10016_ _15202_/Q _15103_/Q _10015_/B vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__a21oi_2
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_76_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__A1 _07732_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12069__B1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__inv_2
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07812__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__B_N _15035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__B _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14755_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14755_/Y sky130_fd_sc_hd__inv_2
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11967_ _11968_/A _11968_/B vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__nor2_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13706_ _13706_/A _13829_/A vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__xor2_1
X_10918_ _11121_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10918_/X sky130_fd_sc_hd__xor2_4
X_14686_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14686_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11898_ _11898_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11899_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13637_ _08750_/A _08750_/B _13636_/B _13636_/A vssd1 vssd1 vccd1 vccd1 _13638_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10849_ _10848_/A _10848_/B _10159_/B vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater545_A _10806_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _13564_/A _13566_/X _13564_/B _13570_/A _13567_/X vssd1 vssd1 vccd1 vccd1
+ _13571_/A sky130_fd_sc_hd__o311a_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15687__D _15687_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A1 _07799_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12792__A1 _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ _15568_/CLK _15307_/D _14359_/Y vssd1 vssd1 vccd1 vccd1 _15307_/Q sky130_fd_sc_hd__dfrtp_1
X_12519_ _14953_/Q _12518_/Y _12517_/A vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__a21o_1
XFILLER_146_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater712_A _15708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ _13499_/A _13499_/B _13584_/A vssd1 vssd1 vccd1 vccd1 _13500_/B sky130_fd_sc_hd__or3_1
X_15238_ _15460_/CLK _15238_/D _14287_/Y vssd1 vssd1 vccd1 vccd1 _15238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_195_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput504 output504/A vssd1 vssd1 vccd1 vccd1 y_r_6[15] sky130_fd_sc_hd__buf_2
XFILLER_160_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput515 _15817_/X vssd1 vssd1 vccd1 vccd1 y_r_7[0] sky130_fd_sc_hd__buf_2
Xoutput526 output526/A vssd1 vssd1 vccd1 vccd1 y_r_7[4] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_29_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15170_/CLK _15169_/D _14213_/Y vssd1 vssd1 vccd1 vccd1 _15169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07991_ _11458_/A _08005_/B _08006_/B vssd1 vssd1 vccd1 vccd1 _07991_/X sky130_fd_sc_hd__or3_1
XFILLER_141_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_119_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09730_ _15096_/Q _15063_/Q vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__or2b_1
XFILLER_171_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10338__B_N _15129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09659_/X _09663_/C vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__and2b_1
XFILLER_67_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08612_ _08728_/B _12945_/A vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__or2_1
XFILLER_54_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09592_ _09590_/X _09597_/B vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07722__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11807__A0 _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ _14912_/Q vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ _14906_/Q vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__buf_6
XFILLER_24_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07425_ _07425_/A vssd1 vssd1 vccd1 vccd1 _15551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07958__A _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 _15416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09026_ _13612_/A _09026_/B vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11199__B _15029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09928_ _15227_/Q _15194_/Q vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__or2b_1
XANTENNA__12104__A _12451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _09859_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _15755_/D sky130_fd_sc_hd__xor2_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07714__A1 _07714_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12870_ _12870_/A _12949_/A vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input126_A x_i_7[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07632__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A _11821_/B _11821_/C vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11662__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14540_/Y sky130_fd_sc_hd__inv_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11832_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__xnor2_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09132__B _15491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10703_ _15281_/Q _15182_/Q vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__and2b_1
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14471_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14471_/Y sky130_fd_sc_hd__inv_2
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11538_/A _11612_/A _11827_/B vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input91_A x_i_5[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ _13422_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__or2_1
XFILLER_197_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10634_ _10634_/A _10634_/B vssd1 vssd1 vccd1 vccd1 _15037_/D sky130_fd_sc_hd__nor2_2
XFILLER_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ _13422_/A _13366_/A _13352_/A vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__a21o_1
X_10565_ _10565_/A _10565_/B _10616_/A vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__and3_1
XFILLER_154_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15300__D _15300_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12304_ _12304_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13284_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__a21o_1
X_10496_ _10496_/A _10496_/B _10592_/A vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__and3_1
X_15023_ _15220_/CLK _15023_/D _14060_/Y vssd1 vssd1 vccd1 vccd1 _15023_/Q sky130_fd_sc_hd__dfrtp_1
X_12235_ _12236_/A _12236_/B _12236_/C vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__o21a_1
XFILLER_194_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07402__A0 _15566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__B _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__nor2_1
XFILLER_151_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11117_ _11117_/A _11117_/B vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12097_ _12096_/B _12096_/C _15735_/Q vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__a21o_1
XFILLER_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11048_ _14928_/Q _14994_/Q vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output512_A _11189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 x_i_0[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12668__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14807_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14807_/Y sky130_fd_sc_hd__inv_2
X_15787_ _15790_/CLK _15787_/D _14867_/Y vssd1 vssd1 vccd1 vccd1 _15787_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _12999_/A _13201_/A _13012_/A vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__or3b_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__A0 _15529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ _14741_/A vssd1 vssd1 vccd1 vccd1 _14738_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14669_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14669_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater927_A input179/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08190_ _08190_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput301 output301/A vssd1 vssd1 vccd1 vccd1 y_i_2[16] sky130_fd_sc_hd__buf_2
XFILLER_173_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput312 _15670_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[10] sky130_fd_sc_hd__buf_2
Xoutput323 output323/A vssd1 vssd1 vccd1 vccd1 y_i_3[5] sky130_fd_sc_hd__buf_2
XFILLER_160_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput334 output334/A vssd1 vssd1 vccd1 vccd1 y_i_4[15] sky130_fd_sc_hd__buf_2
XANTENNA__14404__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput345 _15811_/X vssd1 vssd1 vccd1 vccd1 y_i_5[0] sky130_fd_sc_hd__buf_2
XFILLER_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput356 output356/A vssd1 vssd1 vccd1 vccd1 y_i_5[4] sky130_fd_sc_hd__buf_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput367 output367/A vssd1 vssd1 vccd1 vccd1 y_i_6[14] sky130_fd_sc_hd__buf_2
Xoutput378 _11121_/Y vssd1 vssd1 vccd1 vccd1 y_i_6[9] sky130_fd_sc_hd__buf_2
XFILLER_113_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput389 _15695_/Q vssd1 vssd1 vccd1 vccd1 y_i_7[3] sky130_fd_sc_hd__buf_2
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07974_ _11020_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__and2_1
XFILLER_19_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09713_ _09832_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _15715_/D sky130_fd_sc_hd__xnor2_1
XFILLER_45_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12859__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07960__B _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _09642_/A _09642_/B _09643_/X vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__a21o_1
XFILLER_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10785__A_N _15788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ _15436_/Q _15420_/Q vssd1 vssd1 vccd1 vccd1 _09575_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _08526_/A _08526_/B vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_815 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__inv_2
XFILLER_211_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07408_ _15563_/Q _07408_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08388_ _08410_/B _08388_/B vssd1 vssd1 vccd1 vccd1 _08412_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07632__A0 _15449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ _15164_/Q _15131_/Q vssd1 vssd1 vccd1 vccd1 _10351_/B sky130_fd_sc_hd__and2b_1
XFILLER_136_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _15372_/Q _15356_/Q vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__xnor2_2
XFILLER_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11938__A _12415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _10281_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _15772_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10842__A _10842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14314__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12020_ _15734_/Q _12025_/B vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__xnor2_2
XFILLER_133_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input243_A x_r_7[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__B _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13971_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13971_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15710_ _15777_/CLK _15710_/D _14786_/Y vssd1 vssd1 vccd1 vccd1 _15710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ _13016_/A _13016_/B vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _15705_/CLK _15641_/D _14713_/Y vssd1 vssd1 vccd1 vccd1 _15641_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12853_ _13390_/A _13319_/A vssd1 vssd1 vccd1 vccd1 _12854_/C sky130_fd_sc_hd__xor2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _12238_/A _12122_/A _11803_/C vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__a21oi_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15572_/CLK _15572_/D _14639_/Y vssd1 vssd1 vccd1 vccd1 _15572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_203_922 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12784_ _13046_/A _13220_/A _12784_/C vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__and3_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14523_/Y sky130_fd_sc_hd__inv_2
X_11735_ _12254_/A _12144_/A vssd1 vssd1 vccd1 vccd1 _12071_/B sky130_fd_sc_hd__xor2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14454_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14454_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11666_ _11797_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13405_ _13347_/A _13570_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13406_/B sky130_fd_sc_hd__o21ai_2
XFILLER_70_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ _15263_/Q _15296_/Q vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__and2_1
X_14385_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14385_/Y sky130_fd_sc_hd__inv_2
X_11597_ _11898_/A _12055_/A vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13336_ _13381_/B _13337_/B vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11090__A_N _14935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ _15261_/Q _15294_/Q vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__or2b_1
XANTENNA_output462_A output462/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13267_ _13268_/A _13268_/B vssd1 vssd1 vccd1 vccd1 _13308_/B sky130_fd_sc_hd__and2_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14224__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _10478_/A _10478_/B _10351_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__a21o_1
X_15006_ _15008_/CLK _15006_/D _14042_/Y vssd1 vssd1 vccd1 vccd1 _15006_/Q sky130_fd_sc_hd__dfrtp_1
X_12218_ _12468_/A _12218_/B vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__xor2_4
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08222__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13198_ _13197_/A _13197_/B _13197_/C vssd1 vssd1 vccd1 vccd1 _13274_/A sky130_fd_sc_hd__a21o_1
XFILLER_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12149_ _12149_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater804 _15586_/Q vssd1 vssd1 vccd1 vccd1 output429/A sky130_fd_sc_hd__clkbuf_2
Xrepeater815 _15382_/Q vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__buf_2
Xrepeater826 input89/X vssd1 vssd1 vccd1 vccd1 _07447_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater837 input75/X vssd1 vssd1 vccd1 vccd1 _07604_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater848 input60/X vssd1 vssd1 vccd1 vccd1 _07439_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater877_A input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater859 input46/X vssd1 vssd1 vccd1 vccd1 _07565_/A1 sky130_fd_sc_hd__clkbuf_2
X_07690_ _07690_/A vssd1 vssd1 vccd1 vccd1 _15421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09360_ _15400_/Q _15384_/Q vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__and2b_1
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ _08303_/X _08309_/X _08342_/A _08280_/Y _08310_/Y vssd1 vssd1 vccd1 vccd1
+ _08311_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09291_ _09285_/Y _09289_/B _09287_/B vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10927__A _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13303__A _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07862__A0 _15336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08173_ _08174_/B _08174_/C _08174_/A vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10676__B_N _15277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14134__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08132__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13973__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07957_ _07957_/A vssd1 vssd1 vccd1 vccd1 _07957_/X sky130_fd_sc_hd__buf_6
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08786__B _15322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _15323_/Q _07888_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _15561_/Q _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09631_/C sky130_fd_sc_hd__a21o_1
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _15434_/Q _15418_/Q vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__xnor2_2
XFILLER_43_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A _08509_/B vssd1 vssd1 vccd1 vccd1 _08509_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14954__D _14954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10837__A _10837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14309__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11520_ _15808_/Q vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__buf_4
XFILLER_62_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11451_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input193_A x_r_3[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ _10402_/A _10402_/B vssd1 vssd1 vccd1 vccd1 _14944_/D sky130_fd_sc_hd__nor2_1
XFILLER_183_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14170_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14170_/Y sky130_fd_sc_hd__inv_2
X_11382_ _11382_/A _11382_/B vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__xor2_4
XFILLER_194_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15785__D _15785_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11668__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13124_/C sky130_fd_sc_hd__xnor2_1
X_10333_ _15128_/Q _15161_/Q vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14044__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _12877_/B _13052_/B vssd1 vssd1 vccd1 vccd1 _13057_/C sky130_fd_sc_hd__and2b_1
XANTENNA_input54_A x_i_3[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10264_ _15081_/Q _15246_/Q vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__or2b_1
XFILLER_79_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12003_ _11917_/A _11917_/B _12002_/X vssd1 vssd1 vccd1 vccd1 _12064_/B sky130_fd_sc_hd__a21oi_1
X_10195_ _15071_/Q _15236_/Q vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12905_ _12906_/A _12906_/B _12906_/C vssd1 vssd1 vccd1 vccd1 _12985_/C sky130_fd_sc_hd__a21o_1
XFILLER_189_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13885_ _13885_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _15058_/D sky130_fd_sc_hd__xnor2_1
XFILLER_59_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output308_A _10905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1059 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15624_ _15741_/CLK _15624_/D _14695_/Y vssd1 vssd1 vccd1 vccd1 _15624_/Q sky130_fd_sc_hd__dfrtp_2
X_12836_ _12836_/A _12836_/B _12836_/C vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__nand3_1
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07820__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_932 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09601__A _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15555_ _15576_/CLK _15555_/D _14622_/Y vssd1 vssd1 vccd1 vccd1 _15555_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _13669_/A _13646_/B vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__nand2_2
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14219__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14506_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11718_ _12378_/B _11719_/B vssd1 vssd1 vccd1 vccd1 _11718_/X sky130_fd_sc_hd__or2_1
XFILLER_14_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15486_ _15508_/CLK _15486_/D _14549_/Y vssd1 vssd1 vccd1 vccd1 _15486_/Q sky130_fd_sc_hd__dfrtp_1
X_12698_ _12699_/A _13528_/B vssd1 vssd1 vccd1 vccd1 _15627_/D sky130_fd_sc_hd__xnor2_1
XFILLER_174_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14437_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14437_/Y sky130_fd_sc_hd__inv_2
X_11649_ _12369_/A _12369_/B _12369_/C vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__nand3b_2
Xinput11 x_i_0[2] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput22 x_i_1[12] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
Xinput33 x_i_1[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 x_i_2[3] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14368_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14368_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput55 x_i_3[13] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
Xinput66 x_i_3[9] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput77 x_i_4[4] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15695__D _15695_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput88 x_i_5[14] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_4
X_13319_ _13319_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13340_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput99 x_i_6[0] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14299_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14299_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14889__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ _08859_/Y _15447_/Q _08857_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater601 _10669_/Y vssd1 vssd1 vccd1 vccd1 _15044_/D sky130_fd_sc_hd__clkbuf_2
X_07811_ _07811_/A vssd1 vssd1 vccd1 vccd1 _15362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater612 _11046_/Y vssd1 vssd1 vccd1 vccd1 repeater612/X sky130_fd_sc_hd__buf_2
X_08791_ _13888_/A _08788_/B _08790_/X vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater623 _11359_/Y vssd1 vssd1 vccd1 vccd1 output441/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater634 _11253_/Y vssd1 vssd1 vccd1 vccd1 output473/A sky130_fd_sc_hd__clkbuf_2
Xrepeater645 _10723_/Y vssd1 vssd1 vccd1 vccd1 output404/A sky130_fd_sc_hd__clkbuf_2
X_07742_ _15395_/Q _07742_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__mux2_1
Xrepeater656 _14841_/A vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__buf_6
XFILLER_38_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater667 _14737_/A vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__clkbuf_4
Xrepeater678 _14526_/A vssd1 vssd1 vccd1 vccd1 _14540_/A sky130_fd_sc_hd__buf_6
Xrepeater689 _14176_/A vssd1 vssd1 vccd1 vccd1 _14178_/A sky130_fd_sc_hd__buf_6
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07673_ _15429_/Q input243/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ _09414_/B _09412_/B vssd1 vssd1 vccd1 vccd1 _15268_/D sky130_fd_sc_hd__nor2_1
XFILLER_198_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07730__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11760__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__or2_1
XFILLER_178_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14129__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _15398_/Q _09275_/A vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__or2b_1
XFILLER_21_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08225_ _11842_/C _08243_/A _08225_/C vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__or3_1
XFILLER_194_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13968__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08156_ _08192_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08174_/C sky130_fd_sc_hd__and2_1
XFILLER_165_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08087_ _08290_/B _08087_/B vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_898 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14799__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14949__D _14949_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _15368_/Q _15352_/Q vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__xnor2_2
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1007 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _10950_/A _10950_/B _11137_/A vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__a21oi_2
XFILLER_112_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11951__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _13669_/A _13648_/A _13669_/B vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input206_A x_r_4[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882_ _10881_/A _10881_/C _11111_/A vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07640__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12619_/X _12618_/B _12620_/X vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__o21ai_1
XFILLER_73_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09421__A _15529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14039__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ _15341_/CLK _15340_/D _14394_/Y vssd1 vssd1 vccd1 vccd1 _15340_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_157_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12552_ _12549_/A _12550_/A _12549_/B _12551_/X vssd1 vssd1 vccd1 vccd1 _12553_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08037__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11503_ _11503_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _15578_/D sky130_fd_sc_hd__xnor2_1
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15271_ _15399_/CLK _15271_/D _14322_/Y vssd1 vssd1 vccd1 vccd1 _15271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12483_ _12484_/B _12484_/C _12484_/A vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clk/A sky130_fd_sc_hd__clkbuf_8
X_14222_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__inv_2
X_11434_ _11434_/A _08047_/A vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14153_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14153_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15754_/CLK sky130_fd_sc_hd__clkbuf_16
X_11365_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11365_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_180_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _13438_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _13105_/B sky130_fd_sc_hd__or2_1
X_10316_ _10451_/A _10316_/B vssd1 vssd1 vccd1 vccd1 _15780_/D sky130_fd_sc_hd__xnor2_4
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14084_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14084_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11296_ _11296_/A _11296_/B vssd1 vssd1 vccd1 vccd1 _11296_/X sky130_fd_sc_hd__xor2_4
XFILLER_65_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13035_/A _13102_/C vssd1 vssd1 vccd1 vccd1 _13036_/B sky130_fd_sc_hd__xor2_1
XFILLER_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ _11408_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _15767_/D sky130_fd_sc_hd__xor2_1
XANTENNA__14502__A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _10178_/A _10178_/B vssd1 vssd1 vccd1 vccd1 _15806_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08500__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output425_A output425/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14986_ _15347_/CLK _14986_/D _14020_/Y vssd1 vssd1 vccd1 vccd1 _14986_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13937_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13937_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater575_A _11332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ _13868_/A _13868_/B vssd1 vssd1 vccd1 vccd1 _13869_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ _15052_/Q _12818_/B _12818_/C vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__a21oi_1
X_15607_ _15705_/CLK _15607_/D _14677_/Y vssd1 vssd1 vccd1 vccd1 _15607_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater742_A repeater743/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ _13871_/B _14985_/Q vssd1 vssd1 vccd1 vccd1 _13799_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_773 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15539_/CLK _15538_/D _14604_/Y vssd1 vssd1 vccd1 vccd1 _15538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15469_ _15472_/CLK _15469_/D _14531_/Y vssd1 vssd1 vccd1 vccd1 _15469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08010_ _11658_/A vssd1 vssd1 vccd1 vccd1 _08010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12169__A2 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11101__A _14936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09961_ _15232_/Q vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08912_ _08968_/A _15457_/Q vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__or2b_1
XFILLER_170_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _15190_/Q _15223_/Q vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__or2_1
XANTENNA__14412__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08842_/Y _15331_/Q _08838_/B vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__a21oi_1
XFILLER_170_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08774_ _15337_/Q _15321_/Q vssd1 vssd1 vccd1 vccd1 _08775_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07725_ _07725_/A vssd1 vssd1 vccd1 vccd1 _15404_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07656_ _07656_/A vssd1 vssd1 vccd1 vccd1 _15438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07587_ _15471_/Q input68/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09326_ _15408_/Q _15392_/Q vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__or2b_1
XFILLER_181_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ _09257_/A vssd1 vssd1 vccd1 vccd1 _15245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _08231_/A _08231_/B _08207_/Y vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__a21oi_1
XFILLER_182_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ _09188_/A _09188_/B vssd1 vssd1 vccd1 vccd1 _09189_/C sky130_fd_sc_hd__nor2_1
XFILLER_181_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__xor2_1
XFILLER_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12107__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11150_ _15744_/Q _15022_/Q vssd1 vssd1 vccd1 vccd1 _11150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _10809_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10103_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10591__B2 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11081_ _14933_/Q _14999_/Q vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input156_A x_r_1[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14322__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput201 x_r_4[15] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput212 x_r_5[10] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__clkbuf_2
X_10032_ _15206_/Q _15107_/Q vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput223 x_r_5[6] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__clkbuf_2
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 x_r_6[1] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_4
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 x_r_7[11] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__clkbuf_2
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput256 x_r_7[7] vssd1 vssd1 vccd1 vccd1 input256/X sky130_fd_sc_hd__clkbuf_2
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14841_/A vssd1 vssd1 vccd1 vccd1 _14840_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09135__B _15492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A x_i_0[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14771_/Y sky130_fd_sc_hd__inv_2
X_11983_ _11983_/A _11983_/B vssd1 vssd1 vccd1 vccd1 _12439_/B sky130_fd_sc_hd__xnor2_4
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13722_ _13722_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__nand2_1
X_10934_ _10934_/A vssd1 vssd1 vccd1 vccd1 _10934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13653_ _13813_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__xnor2_4
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10865_ _14956_/Q _14890_/Q vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__nand2_1
X_12604_ _12604_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _15687_/D sky130_fd_sc_hd__xnor2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13584_ _13584_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13585_/B sky130_fd_sc_hd__or2b_1
XFILLER_169_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10796_ _10795_/A _10795_/B _11296_/A vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__a21oi_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15712_/CLK _15323_/D _14376_/Y vssd1 vssd1 vccd1 vccd1 _15323_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _15729_/Q _12534_/B _12529_/B _12530_/X _12531_/X vssd1 vssd1 vccd1 vccd1
+ _12536_/B sky130_fd_sc_hd__a221o_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15254_ _15527_/CLK _15254_/D _14304_/Y vssd1 vssd1 vccd1 vccd1 _15254_/Q sky130_fd_sc_hd__dfrtp_1
X_12466_ _12466_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12468_/C sky130_fd_sc_hd__or2b_1
XANTENNA_output375_A output375/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14205_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _15080_/Q _15245_/Q _11416_/B vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__a21o_1
XFILLER_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15185_ _15202_/CLK _15185_/D _14230_/Y vssd1 vssd1 vccd1 vccd1 _15185_/Q sky130_fd_sc_hd__dfrtp_4
X_12397_ _12398_/A _12398_/B _12588_/A vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__o21a_1
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _11348_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__xor2_2
XFILLER_158_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14067_/Y sky130_fd_sc_hd__inv_2
X_11279_ _15717_/Q _11278_/Y _11277_/B vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14232__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _13020_/A _13018_/B _13020_/B vssd1 vssd1 vccd1 vccd1 _13018_/X sky130_fd_sc_hd__or3_1
XANTENNA_repeater692_A _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13790__B _13790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater957_A input139/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ _15133_/CLK _14969_/D _14002_/Y vssd1 vssd1 vccd1 vccd1 _14969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11591__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ _15509_/Q _07510_/A1 _07538_/S vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__mux2_1
X_08490_ _08486_/A _08486_/B _08548_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08506_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_63_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07441_ _15543_/Q _07441_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07442_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09111_ _15503_/Q _15487_/Q vssd1 vssd1 vccd1 vccd1 _09254_/A sky130_fd_sc_hd__or2b_1
XFILLER_176_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14407__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _15361_/Q _15377_/Q vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13311__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13030__B _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09944_ _15230_/Q _15197_/Q vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__or2b_1
XANTENNA__10670__A _15276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14142__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07455__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08140__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09875_ _09875_/A _09875_/B _09973_/A vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__and3_1
XANTENNA_input9_A x_i_0[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13981__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08825_/A _08825_/B _13905_/A vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__a21o_1
XFILLER_100_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _15660_/D sky130_fd_sc_hd__nand2_2
XFILLER_72_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _15412_/Q _07708_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__mux2_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ _08688_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__xor2_1
XFILLER_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07639_/A vssd1 vssd1 vccd1 vccd1 _15446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ _15272_/Q _15173_/Q vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__or2_1
XFILLER_167_710 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09309_ _09302_/Y _09307_/B _09304_/B vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__o21ai_1
XFILLER_10_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14962__D _14962_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10581_ _15265_/Q _10580_/Y _10579_/B vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__a21oi_1
XFILLER_142_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14317__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12320_ _12322_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _12569_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_640 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11202_ _15750_/Q _11201_/Y _11197_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__a21o_2
X_12182_ _12180_/Y _12182_/B vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13875__B _15318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15793__D _15793_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11133_ _11131_/A _11131_/B _11132_/X vssd1 vssd1 vccd1 vccd1 _11134_/B sky130_fd_sc_hd__a21o_2
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10580__A _15298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14052__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09146__A _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ _11064_/A _11339_/A vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__nand2_1
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _14971_/D sky130_fd_sc_hd__nor2_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _14827_/A vssd1 vssd1 vccd1 vccd1 _14823_/Y sky130_fd_sc_hd__inv_2
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__C _11842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ _11966_/A _11966_/B vssd1 vssd1 vccd1 vccd1 _11968_/B sky130_fd_sc_hd__xnor2_1
X_14754_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14754_/Y sky130_fd_sc_hd__inv_2
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ _14962_/Q _10916_/Y _10912_/B vssd1 vssd1 vccd1 vccd1 _10919_/B sky130_fd_sc_hd__a21o_2
XFILLER_44_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13705_ _14977_/Q _13830_/B vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07496__A1 _07496_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14685_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14685_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11897_ _11898_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__and2_1
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13636_ _13636_/A _13636_/B vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__and2_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10848_ _10848_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _14916_/D sky130_fd_sc_hd__xor2_2
XFILLER_44_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output492_A _15614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13567_ _15767_/Q _13567_/B vssd1 vssd1 vccd1 vccd1 _13567_/X sky130_fd_sc_hd__or2_1
X_10779_ _10779_/A _10779_/B _11292_/A vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__and3_1
XFILLER_201_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14227__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12518_ _12620_/B vssd1 vssd1 vccd1 vccd1 _12518_/Y sky130_fd_sc_hd__inv_2
X_15306_ _15391_/CLK _15306_/D _14358_/Y vssd1 vssd1 vccd1 vccd1 _15306_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__A _11842_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13498_ _13499_/A _13499_/B _13584_/A vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__o21ai_1
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12449_ _12449_/A vssd1 vssd1 vccd1 vccd1 _15652_/D sky130_fd_sc_hd__clkbuf_1
X_15237_ _15477_/CLK _15237_/D _14286_/Y vssd1 vssd1 vccd1 vccd1 _15237_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater705_A _07575_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput505 _11247_/Y vssd1 vssd1 vccd1 vccd1 y_r_6[16] sky130_fd_sc_hd__buf_2
XFILLER_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput516 _15636_/Q vssd1 vssd1 vccd1 vccd1 y_r_7[10] sky130_fd_sc_hd__buf_2
Xoutput527 output527/A vssd1 vssd1 vccd1 vccd1 y_r_7[5] sky130_fd_sc_hd__buf_2
X_15168_ _15775_/CLK _15168_/D _14212_/Y vssd1 vssd1 vccd1 vccd1 _15168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08879__B _15451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__buf_12
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07420__A1 _07420_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _07990_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _08006_/B sky130_fd_sc_hd__xor2_1
XFILLER_140_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15099_ _15375_/CLK _15099_/D _14140_/Y vssd1 vssd1 vccd1 vccd1 _15099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15208__D _15208_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ _09659_/B _09659_/C _09659_/A vssd1 vssd1 vccd1 vccd1 _09663_/C sky130_fd_sc_hd__a21o_1
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08611_ _12708_/A _12871_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _08611_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09591_ _09590_/A _09590_/B _09795_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08542_ _08546_/B _08542_/B vssd1 vssd1 vccd1 vccd1 _08566_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08473_ _14908_/Q vssd1 vssd1 vccd1 vccd1 _12803_/A sky130_fd_sc_hd__buf_6
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07424_ _15551_/Q input52/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10665__A _15275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14137__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08135__A _08223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ _13612_/A _09026_/B vssd1 vssd1 vccd1 vccd1 _15111_/D sky130_fd_sc_hd__xor2_1
XFILLER_156_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13976__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13695__B _13827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12315__A_N _12291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _09987_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09858_ _09857_/A _09857_/B _09743_/B vssd1 vssd1 vccd1 vccd1 _09859_/B sky130_fd_sc_hd__a21o_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14600__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11943__B _11950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _15343_/Q _15327_/Q vssd1 vssd1 vccd1 vccd1 _08818_/A sky130_fd_sc_hd__or2b_1
XFILLER_85_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09789_ _15436_/Q _15420_/Q _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__o21a_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11821_/A _11821_/B _11821_/C vssd1 vssd1 vccd1 vccd1 _11904_/A sky130_fd_sc_hd__a21o_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09413__B _15511_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A x_i_7[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11749_/X _11859_/A vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__and2b_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08029__B _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_80_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15790_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _15280_/Q _15181_/Q vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14470_/Y sky130_fd_sc_hd__inv_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11685_/A sky130_fd_sc_hd__inv_2
XFILLER_14_579 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10582__B_N _15299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ _13422_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13470_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10633_ _10633_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__and2_1
XANTENNA__14047__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_702 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _13352_/A _13422_/A vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input84_A x_i_5[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _10564_/A _10572_/A vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _15739_/Q vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__inv_2
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13283_ _13287_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__xnor2_2
XFILLER_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10495_ _10493_/Y _10495_/B vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ _15444_/CLK _15022_/D _14058_/Y vssd1 vssd1 vccd1 vccd1 _15022_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12236_/C sky130_fd_sc_hd__or2_1
XFILLER_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07402__A1 input126/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _12231_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__xor2_1
XFILLER_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _10891_/Y _11115_/B _10893_/B vssd1 vssd1 vccd1 vccd1 _11117_/B sky130_fd_sc_hd__o21ai_4
XFILLER_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12096_ _15735_/Q _12096_/B _12096_/C vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__and3_1
XFILLER_150_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_890 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output338_A _11308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _14928_/Q _14994_/Q vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__or2_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14510__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 x_i_0[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output505_A _11247_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14806_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15786_ _15790_/CLK _15786_/D _14866_/Y vssd1 vssd1 vccd1 vccd1 _15786_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _13203_/A vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__clkinv_2
XFILLER_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__A1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14737_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14737_/Y sky130_fd_sc_hd__inv_2
X_11949_ _15733_/Q vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__clkinv_2
XANTENNA_repeater655_A _07957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 _15689_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _14681_/A vssd1 vssd1 vccd1 vccd1 _14668_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15698__D _15698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater822_A input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ _13618_/B _13618_/C _13618_/A vssd1 vssd1 vccd1 vccd1 _13620_/B sky130_fd_sc_hd__o21a_1
X_14599_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14599_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput302 output302/A vssd1 vssd1 vccd1 vccd1 y_i_2[1] sky130_fd_sc_hd__buf_2
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput313 output313/A vssd1 vssd1 vccd1 vccd1 y_i_3[11] sky130_fd_sc_hd__buf_2
Xoutput324 _15666_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[6] sky130_fd_sc_hd__buf_2
XFILLER_142_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput335 _11352_/Y vssd1 vssd1 vccd1 vccd1 y_i_4[16] sky130_fd_sc_hd__buf_2
Xoutput346 _15686_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[10] sky130_fd_sc_hd__buf_2
XFILLER_160_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput357 _15681_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[5] sky130_fd_sc_hd__buf_2
XFILLER_142_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput368 output368/A vssd1 vssd1 vccd1 vccd1 y_i_6[15] sky130_fd_sc_hd__buf_2
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput379 _15813_/X vssd1 vssd1 vccd1 vccd1 y_i_7[0] sky130_fd_sc_hd__buf_2
XFILLER_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ _14921_/Q _14987_/Q vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__or2_1
XFILLER_206_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09712_ _09706_/A _09708_/B _09706_/B vssd1 vssd1 vccd1 vccd1 _09713_/B sky130_fd_sc_hd__a21boi_1
XFILLER_68_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14420__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12859__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _15566_/Q _15546_/Q vssd1 vssd1 vccd1 vccd1 _09643_/X sky130_fd_sc_hd__and2b_1
XFILLER_167_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ _09572_/Y _09574_/B vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__nand2b_1
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10379__B _10486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08525_ _08525_/A _08672_/C vssd1 vssd1 vccd1 vccd1 _08526_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_62_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15784_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_60_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ _08600_/A _08619_/A vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__nor2_1
XFILLER_195_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07407_ _07407_/A vssd1 vssd1 vccd1 vccd1 _15564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08387_ _08385_/Y _08447_/B _12627_/A vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07880__A1 input132/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_75_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07632__A1 _07632_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _13605_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _15108_/D sky130_fd_sc_hd__xor2_1
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ _10279_/A _10279_/B _11424_/A vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__a21oi_1
XFILLER_133_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14330__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13970_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input236_A x_r_6[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _12921_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _13016_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15640_ _15771_/CLK _15640_/D _14712_/Y vssd1 vssd1 vccd1 vccd1 _15640_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12851_/Y _12786_/A _12787_/B _12787_/A vssd1 vssd1 vccd1 vccd1 _12867_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _12238_/A _12122_/A _11803_/C vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__and3_1
XFILLER_33_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12970_/A _12871_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _12787_/A sky130_fd_sc_hd__and3b_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15571_/CLK _15571_/D _14638_/Y vssd1 vssd1 vccd1 vccd1 _15571_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_28_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15180_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_1011 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11742_/A _11734_/B _11734_/C vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__or3_1
XFILLER_199_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14522_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _11766_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__nor2_1
X_14453_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14453_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_186_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13404_ _15768_/Q _13572_/A vssd1 vssd1 vccd1 vccd1 _13404_/Y sky130_fd_sc_hd__nand2_1
X_10616_ _10616_/A _10616_/B vssd1 vssd1 vccd1 vccd1 _14999_/D sky130_fd_sc_hd__xor2_1
X_14384_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14384_/Y sky130_fd_sc_hd__inv_2
X_11596_ _11596_/A _11596_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__xor2_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output288_A output288/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13335_ _13335_/A _13393_/A vssd1 vssd1 vccd1 vccd1 _13337_/B sky130_fd_sc_hd__and2_1
X_10547_ _15293_/Q _15260_/Q vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__or2b_1
XFILLER_182_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14505__A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07818__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _13187_/A _13187_/B _13265_/X vssd1 vssd1 vccd1 vccd1 _13268_/B sky130_fd_sc_hd__a21o_1
X_10478_ _10478_/A _10478_/B vssd1 vssd1 vccd1 vccd1 _14900_/D sky130_fd_sc_hd__xor2_1
XANTENNA_output455_A output455/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12217_ _12152_/A _12215_/Y _12216_/Y vssd1 vssd1 vccd1 vccd1 _12218_/B sky130_fd_sc_hd__a21o_1
X_15005_ _15008_/CLK _15005_/D _14041_/Y vssd1 vssd1 vccd1 vccd1 _15005_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_974 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13197_ _13197_/A _13197_/B _13197_/C vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__and3_1
XFILLER_9_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12148_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__and3_1
XFILLER_150_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater805 _15584_/Q vssd1 vssd1 vccd1 vccd1 output427/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater816 _14862_/A vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__buf_6
XFILLER_42_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ _12079_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12132__A0 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater827 input88/X vssd1 vssd1 vccd1 vccd1 _07449_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__14240__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater838 input74/X vssd1 vssd1 vccd1 vccd1 _07606_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater849 input6/X vssd1 vssd1 vccd1 vccd1 _07616_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07553__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _15774_/CLK _15769_/D _14848_/Y vssd1 vssd1 vccd1 vccd1 _15769_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_44_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15008_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ _08310_/A _08310_/B vssd1 vssd1 vccd1 vccd1 _08310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09290_ _15401_/Q _15385_/Q vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__xnor2_2
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08241_ _08254_/A _08253_/A vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__or2_1
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07862__A1 input204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08172_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__xor2_1
XFILLER_192_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07614__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_919 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14415__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07728__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09228__B _15480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08132__B _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07956_ _11105_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__and2_1
XFILLER_130_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14150__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07887_ _07887_/A vssd1 vssd1 vccd1 vccd1 _15324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _15541_/Q vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__inv_2
XFILLER_16_619 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _09781_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _15172_/D sky130_fd_sc_hd__xor2_1
XFILLER_15_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15406_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08508_ _08503_/B _08508_/B vssd1 vssd1 vccd1 vccd1 _08528_/A sky130_fd_sc_hd__and2b_1
XFILLER_145_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09488_ _15540_/Q _15524_/Q vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__or2_1
XFILLER_93_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08439_ _13203_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08458_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15131__D _15131_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _11450_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__xnor2_1
X_10401_ _10400_/B _10400_/C _10400_/A vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14970__D _14970_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11379_/A _11379_/B _11380_/X vssd1 vssd1 vccd1 vccd1 _11382_/B sky130_fd_sc_hd__a21o_1
XFILLER_194_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14325__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_671 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input186_A x_r_3[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13144_/B _13120_/B vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07638__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _15128_/Q _15161_/Q vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__or2_1
XANTENNA__11668__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ _13054_/A _13054_/B vssd1 vssd1 vccd1 vccd1 _13051_/Y sky130_fd_sc_hd__nand2_1
X_10263_ _10263_/A vssd1 vssd1 vccd1 vccd1 _15769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _11916_/B _12002_/B vssd1 vssd1 vccd1 vccd1 _12002_/X sky130_fd_sc_hd__and2b_1
XFILLER_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A x_i_2[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10194_ _15071_/Q _15236_/Q vssd1 vssd1 vccd1 vccd1 _10194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14060__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13953_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12921_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _12906_/C sky130_fd_sc_hd__xnor2_1
XFILLER_98_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08993__A _15369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A0 _15494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13884_ _08773_/Y _13883_/B _08775_/B vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__o21ai_2
XFILLER_35_939 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15623_ _15717_/CLK _15623_/D _14694_/Y vssd1 vssd1 vccd1 vccd1 _15623_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_991 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12836_/A _12836_/B _12836_/C vssd1 vssd1 vccd1 vccd1 _12835_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15400_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15569_/CLK _15554_/D _14620_/Y vssd1 vssd1 vccd1 vccd1 _15554_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12766_ _12777_/A _12777_/B _12775_/A vssd1 vssd1 vccd1 vccd1 _13646_/B sky130_fd_sc_hd__nand3_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14505_/Y sky130_fd_sc_hd__inv_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11727_/A _11717_/B vssd1 vssd1 vccd1 vccd1 _12381_/A sky130_fd_sc_hd__and2_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07844__A1 _07844_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12697_ _12700_/A _13529_/B vssd1 vssd1 vccd1 vccd1 _13528_/B sky130_fd_sc_hd__xnor2_2
X_15485_ _15571_/CLK _15485_/D _14548_/Y vssd1 vssd1 vccd1 vccd1 _15485_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15041__D _15041_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__or2_1
XFILLER_174_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14436_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14436_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput12 x_i_0[3] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
Xinput23 x_i_1[13] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput34 x_i_1[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput45 x_i_2[4] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
X_11579_ _15728_/Q _11581_/B vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__xor2_2
X_14367_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14367_/Y sky130_fd_sc_hd__inv_2
Xinput56 x_i_3[14] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14235__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_811 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 x_i_4[0] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput78 x_i_4[5] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
Xinput89 x_i_5[15] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_2
X_13318_ _13318_/A _13318_/B vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__xnor2_2
XFILLER_192_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14298_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14298_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__or2_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07810_ _15362_/Q input167/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08790_ _15339_/Q _15323_/Q vssd1 vssd1 vccd1 vccd1 _08790_/X sky130_fd_sc_hd__and2b_1
Xrepeater602 _11365_/Y vssd1 vssd1 vccd1 vccd1 output444/A sky130_fd_sc_hd__clkbuf_2
Xrepeater613 _10889_/X vssd1 vssd1 vccd1 vccd1 output306/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater624 _11111_/Y vssd1 vssd1 vccd1 vccd1 output373/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater635 repeater636/X vssd1 vssd1 vccd1 vccd1 output507/A sky130_fd_sc_hd__buf_4
XFILLER_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ _07741_/A vssd1 vssd1 vccd1 vccd1 _15396_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater646 _11353_/Y vssd1 vssd1 vccd1 vccd1 output438/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater657 _14827_/A vssd1 vssd1 vccd1 vccd1 _14841_/A sky130_fd_sc_hd__buf_6
XFILLER_37_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater668 _14737_/A vssd1 vssd1 vccd1 vccd1 _14740_/A sky130_fd_sc_hd__buf_6
XFILLER_203_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater679 _14526_/A vssd1 vssd1 vccd1 vccd1 _14538_/A sky130_fd_sc_hd__buf_6
X_07672_ _07672_/A vssd1 vssd1 vccd1 vccd1 _15430_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09411_ _15525_/Q _09411_/B _09495_/B vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__and3_1
XFILLER_52_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15192_/CLK sky130_fd_sc_hd__clkbuf_16
X_09342_ _15412_/Q _15396_/Q vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__nor2_1
XFILLER_205_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _09271_/A _09271_/B _09272_/X vssd1 vssd1 vccd1 vccd1 _15250_/D sky130_fd_sc_hd__a21o_1
XFILLER_193_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ _11491_/A _08223_/B _08223_/C vssd1 vssd1 vccd1 vccd1 _08225_/C sky130_fd_sc_hd__a21oi_1
XFILLER_20_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08192_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14145__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ _08086_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__xor2_2
XANTENNA__08143__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13984__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07982__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07771__A0 _15381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08988_ _08988_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _15104_/D sky130_fd_sc_hd__nor2_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _07939_/A _10380_/A vssd1 vssd1 vccd1 vccd1 _10014_/A sky130_fd_sc_hd__nor2_1
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09512__A1 _15532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _10950_/A _10950_/B _11137_/A vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__and3_1
XFILLER_44_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09609_ _15442_/Q _15426_/Q vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__and2b_1
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10881_ _10881_/A _11111_/A _10881_/C vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__and3_1
XFILLER_204_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13224__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _14953_/Q _12620_/B vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__or2_1
XANTENNA_input101_A x_i_6[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08318__A _15726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_931 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12551_ _12223_/A _12223_/B _15734_/Q vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07826__A1 input174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11502_ _15727_/Q _12527_/B vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__xnor2_2
XFILLER_145_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ _12482_/A _12213_/A vssd1 vssd1 vccd1 vccd1 _12484_/C sky130_fd_sc_hd__or2b_1
X_15270_ _15399_/CLK _15270_/D _14321_/Y vssd1 vssd1 vccd1 vccd1 _15270_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15796__D _15796_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _08123_/A _08123_/B _11432_/X vssd1 vssd1 vccd1 vccd1 _11463_/A sky130_fd_sc_hd__a21oi_2
XFILLER_172_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14221_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14221_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14055__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__A _15299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09149__A _15563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14152_/Y sky130_fd_sc_hd__inv_2
X_11364_ _11177_/Y _11363_/B _11179_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__08053__A _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10315_ _10307_/Y _10311_/B _10309_/B vssd1 vssd1 vccd1 vccd1 _10316_/B sky130_fd_sc_hd__o21ai_4
XFILLER_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _13438_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__nand2_1
X_14083_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14083_/Y sky130_fd_sc_hd__inv_2
X_11295_ _11294_/A _11294_/B _10786_/B vssd1 vssd1 vccd1 vccd1 _11296_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13034_ _13034_/A _13034_/B vssd1 vssd1 vccd1 vccd1 _13102_/C sky130_fd_sc_hd__xnor2_1
XFILLER_152_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10246_ _15077_/Q _10245_/Y _10241_/B vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11543__D1 _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10177_ _10176_/A _10176_/B _10852_/A vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__a21oi_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output320_A _15662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14985_ _15347_/CLK _14985_/D _14019_/Y vssd1 vssd1 vccd1 vccd1 _14985_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_output418_A _15591_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13936_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07514__A0 _15507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13867_ _13867_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _13868_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13688__C_N _12976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater568_A _11379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15606_ _15770_/CLK _15606_/D _14676_/Y vssd1 vssd1 vccd1 vccd1 _15606_/Q sky130_fd_sc_hd__dfrtp_2
X_12818_ _15052_/Q _12818_/B _12818_/C vssd1 vssd1 vccd1 vccd1 _12820_/A sky130_fd_sc_hd__and3_1
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13798_ _13869_/A vssd1 vssd1 vccd1 vccd1 _13798_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _15539_/CLK _15537_/D _14603_/Y vssd1 vssd1 vccd1 vccd1 _15537_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater735_A _15671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _12800_/A sky130_fd_sc_hd__xor2_1
XFILLER_188_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15468_ _15558_/CLK _15468_/D _14530_/Y vssd1 vssd1 vccd1 vccd1 _15468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14419_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater902_A input219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ _15399_/CLK _15399_/D _14457_/Y vssd1 vssd1 vccd1 vccd1 _15399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11101__B _15002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _14968_/D sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_6_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15558_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08898__A _15471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _15457_/Q _08968_/A vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__or2b_1
XFILLER_174_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09891_ _09891_/A _09896_/A vssd1 vssd1 vccd1 vccd1 _14958_/D sky130_fd_sc_hd__nor2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08842_ _15347_/Q vssd1 vssd1 vccd1 vccd1 _08842_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12213__A _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12629__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _15337_/Q _15321_/Q vssd1 vssd1 vccd1 vccd1 _08773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07724_ _15404_/Q input224/X _07750_/S vssd1 vssd1 vccd1 vccd1 _07725_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_894 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07655_ _15438_/Q input258/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07656_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07586_ _07586_/A vssd1 vssd1 vccd1 vccd1 _15472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1071 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09325_ _15392_/Q _15408_/Q vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__or2b_1
XFILLER_159_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13979__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07808__A1 _07808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09254_/X _09258_/C vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__and2b_1
XFILLER_139_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09187_ _09187_/A _09663_/A vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ _08157_/A _08223_/C _11491_/A vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__B _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _08290_/B _08069_/B vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__nor2_1
XFILLER_175_1056 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14603__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _15136_/Q _15301_/Q vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__or2b_1
XFILLER_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11080_ _11080_/A vssd1 vssd1 vccd1 vccd1 _11080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput202 x_r_4[1] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_4
X_10031_ _15206_/Q _15107_/Q vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__or2_1
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 x_r_5[11] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput224 x_r_5[7] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__clkbuf_2
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input149_A x_r_1[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput235 x_r_6[2] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__clkbuf_1
Xinput246 x_r_7[12] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__clkbuf_2
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput257 x_r_7[8] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__clkbuf_1
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14770_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13293__A1 _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ _11904_/A _11904_/B _11903_/A _11902_/A vssd1 vssd1 vccd1 vccd1 _11983_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07651__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_894 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _13721_/A _13832_/B vssd1 vssd1 vccd1 vccd1 _15700_/D sky130_fd_sc_hd__xor2_1
XFILLER_99_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10933_ _10931_/X _10938_/B vssd1 vssd1 vccd1 vccd1 _10933_/X sky130_fd_sc_hd__and2b_2
XFILLER_16_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10864_ _14956_/Q _14890_/Q vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__nor2_1
X_13652_ _13652_/A _13652_/B vssd1 vssd1 vccd1 vccd1 _13813_/B sky130_fd_sc_hd__xor2_4
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _12601_/A _12601_/B _12602_/X vssd1 vssd1 vccd1 vccd1 _12604_/B sky130_fd_sc_hd__a21oi_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13596__A2 _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10795_ _10795_/A _10795_/B _11296_/A vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__and3_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13584_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _15608_/D sky130_fd_sc_hd__xnor2_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15774_/CLK _15322_/D _14375_/Y vssd1 vssd1 vccd1 vccd1 _15322_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12534_ _15729_/Q _12534_/B vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__or2_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _15561_/CLK _15253_/D _14303_/Y vssd1 vssd1 vccd1 vccd1 _15253_/Q sky130_fd_sc_hd__dfrtp_1
X_12465_ _12601_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _15653_/D sky130_fd_sc_hd__xnor2_1
XFILLER_8_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08224__A1 _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _15737_/D sky130_fd_sc_hd__nor2_2
XANTENNA_output270_A output270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12396_ _12396_/A _12395_/Y vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__or2b_1
X_15184_ _15184_/CLK _15184_/D _14229_/Y vssd1 vssd1 vccd1 vccd1 _15184_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output368_A output368/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ _11346_/A _11346_/B _11084_/B vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__a21o_2
X_14135_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14135_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09972__B2 _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14513__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07826__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11278_ _15783_/Q vssd1 vssd1 vccd1 vccd1 _11278_/Y sky130_fd_sc_hd__inv_2
X_14066_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14066_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10760__B _15784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13017_ _13017_/A _12946_/A vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__or2b_1
X_10229_ _15076_/Q _15241_/Q vssd1 vssd1 vccd1 vccd1 _10230_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12033__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater685_A _14439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14968_ _15428_/CLK _14968_/D _14001_/Y vssd1 vssd1 vccd1 vccd1 _14968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07561__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13919_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater852_A repeater853/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A _15252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14899_ _15729_/CLK _14899_/D _13928_/Y vssd1 vssd1 vccd1 vccd1 _14899_/Q sky130_fd_sc_hd__dfrtp_1
X_07440_ _07440_/A vssd1 vssd1 vccd1 vccd1 _15544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_870 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09110_ _15487_/Q _15503_/Q vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__or2b_1
XFILLER_31_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ _09041_/A vssd1 vssd1 vccd1 vccd1 _15113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14423__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07736__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _15197_/Q _15230_/Q vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__or2b_1
XFILLER_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08421__A _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09874_ _09872_/Y _09874_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__and2b_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08825_ _08825_/A _08825_/B _13905_/A vssd1 vssd1 vccd1 vccd1 _08825_/X sky130_fd_sc_hd__and3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _14938_/Q _13808_/A vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nand2_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07471__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07707_ _07707_/A vssd1 vssd1 vccd1 vccd1 _15413_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10981__B_N _15272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10398__A _10398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08687_ _12680_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _08688_/B sky130_fd_sc_hd__xor2_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _15446_/Q input10/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__mux2_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07569_ _15480_/Q input44/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07570_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ _15405_/Q _15389_/Q vssd1 vssd1 vccd1 vccd1 _09375_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ _15298_/Q vssd1 vssd1 vccd1 vccd1 _10580_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _15241_/D sky130_fd_sc_hd__xor2_2
XFILLER_194_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12252_/C sky130_fd_sc_hd__or2_1
XFILLER_177_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _15028_/Q vssd1 vssd1 vccd1 vccd1 _11201_/Y sky130_fd_sc_hd__inv_2
X_12181_ _12181_/A _12181_/B _12181_/C vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nand3_1
XFILLER_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14333__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A1 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ _14966_/Q _14900_/Q vssd1 vssd1 vccd1 vccd1 _11132_/X sky130_fd_sc_hd__and2_1
XFILLER_107_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_654 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ _14997_/Q _14931_/Q vssd1 vssd1 vccd1 vccd1 _11339_/A sky130_fd_sc_hd__or2b_1
XANTENNA__09146__B _15541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10014_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__and2_1
XFILLER_209_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08985__B _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14827_/A sky130_fd_sc_hd__buf_6
XANTENNA__12069__A2 _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09162__A _15566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14753_/Y sky130_fd_sc_hd__inv_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _11963_/X _11965_/B vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__and2b_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13704_ _13704_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__xnor2_4
X_10916_ _14896_/Q vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__inv_2
X_14684_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14684_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11896_ _11953_/B _11896_/B vssd1 vssd1 vccd1 vccd1 _11898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _13649_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13639_/A sky130_fd_sc_hd__xnor2_2
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ _15146_/Q _10846_/Y _10845_/B vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14508__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ _15767_/Q _13567_/B vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__and2_1
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10778_ _10778_/A _10778_/B vssd1 vssd1 vccd1 vccd1 _11292_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output485_A _15623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ _15592_/CLK _15305_/D _14357_/Y vssd1 vssd1 vccd1 vccd1 _15305_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12737__A_N _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _15658_/D sky130_fd_sc_hd__nor2_1
XFILLER_158_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _13585_/A _13497_/B vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__nand2_1
XFILLER_201_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15236_ _15464_/CLK _15236_/D _14285_/Y vssd1 vssd1 vccd1 vccd1 _15236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12448_ _12464_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12449_/A sky130_fd_sc_hd__and2_1
XFILLER_138_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput506 output506/A vssd1 vssd1 vccd1 vccd1 y_r_6[1] sky130_fd_sc_hd__buf_2
XFILLER_176_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput517 output517/A vssd1 vssd1 vccd1 vccd1 y_r_7[11] sky130_fd_sc_hd__buf_2
X_15167_ _15777_/CLK _15167_/D _14211_/Y vssd1 vssd1 vccd1 vccd1 _15167_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput528 _15632_/Q vssd1 vssd1 vccd1 vccd1 y_r_7[6] sky130_fd_sc_hd__buf_2
X_12379_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12381_/D sky130_fd_sc_hd__inv_2
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14243__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14118_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15098_ _15375_/CLK _15098_/D _14138_/Y vssd1 vssd1 vccd1 vccd1 _15098_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14049_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14049_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ _12630_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _08732_/B sky130_fd_sc_hd__and2_1
X_09590_ _09590_/A _09590_/B _09795_/B vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__and3_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08387__S _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_274 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08541_ _08550_/A _08536_/C _13030_/C vssd1 vssd1 vccd1 vccd1 _08542_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1003 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _12780_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08478_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07423_ _07423_/A vssd1 vssd1 vccd1 vccd1 _15552_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10491__A1 _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14418__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13322__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _13610_/A _09018_/B _09023_/X vssd1 vssd1 vccd1 vccd1 _09026_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10681__A _15277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14153__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08151__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13992__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _09987_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _14963_/D sky130_fd_sc_hd__xor2_2
XFILLER_120_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _15754_/D sky130_fd_sc_hd__xor2_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _15327_/Q _15343_/Q vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__or2b_1
XFILLER_6_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _15159_/D sky130_fd_sc_hd__xnor2_1
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _08722_/Y _08723_/X _08724_/X _08725_/X _08738_/X vssd1 vssd1 vccd1 vccd1
+ _08739_/X sky130_fd_sc_hd__a221o_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15134__D _15134_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11749_/A _11749_/B _11749_/C vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__a21o_1
XFILLER_121_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10701_/A vssd1 vssd1 vccd1 vccd1 _15049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14973__D _14973_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__or2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14328__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13420_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__xor2_1
X_10632_ _10633_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13351_ _13351_/A _13307_/A vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__or2b_1
X_10563_ _15296_/Q _15263_/Q vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__or2b_1
XFILLER_195_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _12302_/A vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__inv_2
XANTENNA_input77_A x_i_4[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10494_ _15253_/Q _15286_/Q vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__nand2_1
X_13282_ _13282_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13567_/B sky130_fd_sc_hd__xnor2_4
XFILLER_5_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11687__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _15444_/CLK _15021_/D _14057_/Y vssd1 vssd1 vccd1 vccd1 _15021_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _12164_/A _12231_/Y _12230_/X _12229_/Y vssd1 vssd1 vccd1 vccd1 _12234_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_170_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14063__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12164_ _12164_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__nand2_1
XFILLER_190_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_123_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12095_ _12428_/A _12223_/A _12455_/C vssd1 vssd1 vccd1 vccd1 _12096_/C sky130_fd_sc_hd__o21ai_1
XFILLER_7_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11046_ _11319_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11046_/Y sky130_fd_sc_hd__xnor2_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13407__A _13576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14805_/Y sky130_fd_sc_hd__inv_2
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _15790_/CLK _15785_/D _14865_/Y vssd1 vssd1 vccd1 vccd1 _15785_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ _13192_/B _12997_/B vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15044__D _15044_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14736_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14736_/Y sky130_fd_sc_hd__inv_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ _11948_/A vssd1 vssd1 vccd1 vccd1 _15584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_206_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _14681_/A vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater550_A _11292_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _12238_/A _12231_/A vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14238__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13618_ _13618_/A _13618_/B _13618_/C vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__nor3_1
XFILLER_38_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__A _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14598_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14598_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _13549_/A _13549_/B vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__and2_1
XFILLER_186_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput303 output303/A vssd1 vssd1 vccd1 vccd1 y_i_2[2] sky130_fd_sc_hd__buf_2
X_15219_ _15444_/CLK _15219_/D _14267_/Y vssd1 vssd1 vccd1 vccd1 _15219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput314 output314/A vssd1 vssd1 vccd1 vccd1 y_i_3[12] sky130_fd_sc_hd__buf_2
XFILLER_127_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput325 output325/A vssd1 vssd1 vccd1 vccd1 y_i_3[7] sky130_fd_sc_hd__buf_2
Xoutput336 output336/A vssd1 vssd1 vccd1 vccd1 y_i_4[1] sky130_fd_sc_hd__buf_2
Xoutput347 _15687_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[11] sky130_fd_sc_hd__buf_2
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09067__A _15494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput358 _15682_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[6] sky130_fd_sc_hd__buf_2
Xoutput369 _11143_/Y vssd1 vssd1 vccd1 vccd1 y_i_6[16] sky130_fd_sc_hd__buf_2
XFILLER_99_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07972_ _14921_/Q _14987_/Q vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__nand2_2
XANTENNA__14701__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ _09709_/Y _09711_/B vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__and2b_1
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _15305_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09573_ _15437_/Q _15421_/Q vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ _08524_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _08672_/C sky130_fd_sc_hd__xor2_1
XFILLER_208_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08455_ _08455_/A _08455_/B _08613_/A vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__or3_1
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14148__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07406_ _15564_/Q input124/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__mux2_1
X_08386_ _08396_/A _12654_/A vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__xor2_1
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13987__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12891__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11964__A1 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A2 _15784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09007_ _13602_/A _09002_/B _09006_/X vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__a21o_1
XFILLER_164_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07396__A1 _07396_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14611__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14968__D _14968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13227__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _12918_/A _13541_/A _12919_/X vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__a21oi_2
XFILLER_76_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input131_A x_r_0[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09424__B _15512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input229_A x_r_6[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ _12970_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11882_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11803_/C sky130_fd_sc_hd__and2_1
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15571_/CLK _15570_/D _14637_/Y vssd1 vssd1 vccd1 vccd1 _15570_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12741_/A _12741_/B _12781_/Y vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__a21bo_1
XFILLER_14_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15799__D _15799_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14526_/A sky130_fd_sc_hd__buf_6
X_11733_ _11733_/A _11705_/A vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__or2b_1
XFILLER_109_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14058__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14452_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14452_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _12122_/A _11977_/A _11663_/C vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__a21oi_1
XFILLER_70_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _13403_/A vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__clkinv_2
XFILLER_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ _15262_/Q _15295_/Q _10614_/B vssd1 vssd1 vccd1 vccd1 _10616_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09073__A1 _15494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14383_/Y sky130_fd_sc_hd__inv_2
X_11595_ _11595_/A _11595_/B _11594_/X vssd1 vssd1 vccd1 vccd1 _11596_/B sky130_fd_sc_hd__or3b_1
XFILLER_168_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _13333_/A _13333_/B _13333_/C vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__o21ai_1
X_10546_ _10546_/A vssd1 vssd1 vccd1 vccd1 _15029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ _13186_/B _13265_/B vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__and2b_1
X_10477_ _15130_/Q _10476_/Y _10475_/B vssd1 vssd1 vccd1 vccd1 _10478_/B sky130_fd_sc_hd__a21o_1
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15170_/CLK _15004_/D _14040_/Y vssd1 vssd1 vccd1 vccd1 _15004_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _12466_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output350_A output350/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _13270_/B _13196_/B vssd1 vssd1 vccd1 vccd1 _13197_/C sky130_fd_sc_hd__nand2_1
XANTENNA_output448_A output448/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15039__D _15039_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _12209_/A _12209_/B vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__xnor2_2
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07834__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater806 _15583_/Q vssd1 vssd1 vccd1 vccd1 output426/A sky130_fd_sc_hd__clkbuf_2
X_12078_ _12079_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__and2_1
Xrepeater817 _07699_/A vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__buf_6
XFILLER_81_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater828 input87/X vssd1 vssd1 vccd1 vccd1 _07451_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater839 input69/X vssd1 vssd1 vccd1 vccd1 _07585_/A1 sky130_fd_sc_hd__buf_4
XANTENNA_repeater598_A _11056_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ _11029_/A _11029_/B vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__nand2_4
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_594 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater765_A _15634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11880__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15768_ _15768_/CLK _15768_/D _14847_/Y vssd1 vssd1 vccd1 vccd1 _15768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14719_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15699_ _15699_/CLK _15699_/D _14774_/Y vssd1 vssd1 vccd1 vccd1 _15699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _11928_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08171_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _08172_/B sky130_fd_sc_hd__xor2_1
XFILLER_119_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11104__B _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12216__A _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09595__B_N _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14431__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07744__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07955_ _14921_/Q _15775_/Q vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__or2_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09244__B _15485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07886_ _15324_/Q _07886_/A1 _07892_/S vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09625_ _09812_/A _09623_/B _09624_/X vssd1 vssd1 vccd1 vccd1 _15184_/D sky130_fd_sc_hd__a21o_1
XFILLER_55_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09556_ _09778_/A _09551_/B _09555_/X vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__a21o_1
XFILLER_110_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ _08552_/A _08552_/B _08506_/X vssd1 vssd1 vccd1 vccd1 _08697_/B sky130_fd_sc_hd__o21ai_1
XFILLER_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09487_ _15540_/Q _15524_/Q vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__nand2_1
XFILLER_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08438_ _15044_/Q vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__buf_6
XFILLER_11_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _08369_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _08395_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14606__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _10400_/A _10400_/B _10400_/C vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__and3_1
XFILLER_109_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11380_ _15754_/Q _15032_/Q vssd1 vssd1 vccd1 vccd1 _11380_/X sky130_fd_sc_hd__and2_1
XFILLER_165_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10461_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _15783_/D sky130_fd_sc_hd__xnor2_2
XFILLER_139_1016 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input179_A x_r_3[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13050_ _13126_/A _13050_/B vssd1 vssd1 vccd1 vccd1 _13059_/A sky130_fd_sc_hd__xor2_2
X_10262_ _10260_/X _10267_/B vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__and2b_1
XFILLER_191_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _12063_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12064_/A sky130_fd_sc_hd__xnor2_1
X_10193_ _15053_/Q _10191_/Y _10197_/B vssd1 vssd1 vccd1 vccd1 _15759_/D sky130_fd_sc_hd__o21a_1
XFILLER_191_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14341__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13952_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13952_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09154__B _15544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09318__B_N _15391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _13016_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__and2_1
XFILLER_98_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13883_ _13883_/A _13883_/B vssd1 vssd1 vccd1 vccd1 _15057_/D sky130_fd_sc_hd__xor2_1
XFILLER_19_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__A1 input106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ _15724_/CLK _15622_/D _14693_/Y vssd1 vssd1 vccd1 vccd1 _15622_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12834_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _12836_/C sky130_fd_sc_hd__xnor2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__B _13572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15553_ _15553_/CLK _15553_/D _14619_/Y vssd1 vssd1 vccd1 vccd1 _15553_/Q sky130_fd_sc_hd__dfrtp_1
X_12765_ _12777_/A _12777_/B _12775_/A vssd1 vssd1 vccd1 vccd1 _13669_/A sky130_fd_sc_hd__a21o_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14504_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14504_/Y sky130_fd_sc_hd__inv_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__A _15029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11716_ _11728_/A _12390_/A vssd1 vssd1 vccd1 vccd1 _11717_/B sky130_fd_sc_hd__nand2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15511_/CLK _15484_/D _14547_/Y vssd1 vssd1 vccd1 vccd1 _15484_/Q sky130_fd_sc_hd__dfrtp_4
X_12696_ _12696_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13529_/B sky130_fd_sc_hd__xnor2_2
XFILLER_203_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output398_A output398/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14435_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14435_/Y sky130_fd_sc_hd__inv_2
X_11647_ _12378_/B _11719_/B vssd1 vssd1 vccd1 vccd1 _12372_/B sky130_fd_sc_hd__xnor2_2
XFILLER_174_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 x_i_0[4] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14516__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 x_i_1[14] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 x_i_2[0] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14366_/Y sky130_fd_sc_hd__inv_2
Xinput46 x_i_2[5] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
X_11578_ _11578_/A _12371_/A vssd1 vssd1 vccd1 vccd1 _11581_/B sky130_fd_sc_hd__xnor2_2
Xinput57 x_i_3[15] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput68 x_i_4[10] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13317_ _13317_/A _13317_/B vssd1 vssd1 vccd1 vccd1 _13318_/B sky130_fd_sc_hd__or2_1
XFILLER_6_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput79 x_i_4[6] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_2
X_10529_ _10600_/A _10524_/B _10528_/X vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__a21o_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14297_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13248_ _13248_/A _13248_/B vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__xor2_4
XFILLER_170_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _13352_/A _15052_/Q vssd1 vssd1 vccd1 vccd1 _13180_/C sky130_fd_sc_hd__nor2_1
XANTENNA__14251__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater603 _11051_/Y vssd1 vssd1 vccd1 vccd1 output274/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater882_A input244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater614 _10748_/Y vssd1 vssd1 vccd1 vccd1 output409/A sky130_fd_sc_hd__clkbuf_2
Xrepeater625 _11036_/Y vssd1 vssd1 vccd1 vccd1 output271/A sky130_fd_sc_hd__clkbuf_2
X_07740_ _15396_/Q _07740_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__mux2_1
Xrepeater636 _11155_/Y vssd1 vssd1 vccd1 vccd1 repeater636/X sky130_fd_sc_hd__buf_2
Xrepeater647 _11105_/Y vssd1 vssd1 vccd1 vccd1 output370/A sky130_fd_sc_hd__clkbuf_2
Xrepeater658 _14787_/A vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__buf_8
XFILLER_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater669 _14709_/A vssd1 vssd1 vccd1 vccd1 _14721_/A sky130_fd_sc_hd__buf_6
XFILLER_37_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07671_ _15430_/Q input250/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07532__A1 _07532_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09410_ _15525_/Q _09411_/B _09495_/B vssd1 vssd1 vccd1 vccd1 _09414_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11220__B_N _15032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09341_ _15412_/Q _15396_/Q vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__and2_1
XFILLER_209_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_89_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15810__A _15810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _15508_/Q _15492_/Q vssd1 vssd1 vccd1 vccd1 _09272_/X sky130_fd_sc_hd__and2b_1
XFILLER_21_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_132_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08223_ _11491_/A _08223_/B _08223_/C vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__and3_1
XFILLER_165_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14426__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _11491_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12592__A1 _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_672 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08085_ _08086_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08272_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08143__B _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__B _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14161__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _08986_/A _08986_/B _13594_/A vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__o21a_1
XFILLER_130_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07771__A1 _07771_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_57_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ _15185_/Q vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__clkinv_2
XFILLER_60_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _07869_/A vssd1 vssd1 vccd1 vccd1 _15333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09608_ _15426_/Q _15442_/Q vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__and2b_1
X_10880_ _14891_/Q _14957_/Q vssd1 vssd1 vccd1 vccd1 _10881_/C sky130_fd_sc_hd__or2b_1
XFILLER_28_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _15414_/Q _15430_/Q vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13224__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _12550_/A _12550_/B vssd1 vssd1 vccd1 vccd1 _15618_/D sky130_fd_sc_hd__xnor2_1
XFILLER_12_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_943 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _12355_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__xor2_2
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14981__D _14981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12481_ _14950_/Q vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__inv_2
XFILLER_138_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14336__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07649__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14220_/Y sky130_fd_sc_hd__inv_2
X_11432_ _08068_/A _11432_/B vssd1 vssd1 vccd1 vccd1 _11432_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12032__B1 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14151_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14151_/Y sky130_fd_sc_hd__inv_2
X_11363_ _11363_/A _11363_/B vssd1 vssd1 vccd1 vccd1 _11363_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_152_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _13162_/B _13102_/B _13102_/C vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__or3_1
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__nand2_2
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14082_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14082_/Y sky130_fd_sc_hd__inv_2
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11294_/X sky130_fd_sc_hd__xor2_1
XFILLER_180_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11695__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ _13116_/B _13033_/B vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__xnor2_1
X_10245_ _15242_/Q vssd1 vssd1 vccd1 vccd1 _10245_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14071__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__C1 _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07384__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10176_ _10176_/A _10176_/B _10852_/A vssd1 vssd1 vccd1 vccd1 _10178_/A sky130_fd_sc_hd__and3_1
XFILLER_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14984_ _15764_/CLK _14984_/D _14017_/Y vssd1 vssd1 vccd1 vccd1 _14984_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13935_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09503__A2 _15512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output313_A output313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07514__A1 _07514_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12957__C _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ _14984_/Q vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__inv_2
XFILLER_35_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _15717_/CLK _15605_/D _14675_/Y vssd1 vssd1 vccd1 vccd1 _15605_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ _12817_/A _12893_/C vssd1 vssd1 vccd1 vccd1 _12818_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13134__B _13558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13797_ _13869_/A _13797_/B vssd1 vssd1 vccd1 vccd1 _15707_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__15052__D _15052_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15536_ _15563_/CLK _15536_/D _14602_/Y vssd1 vssd1 vccd1 vccd1 _15536_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12795_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12749_/B sky130_fd_sc_hd__xor2_1
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ _15467_/CLK _15467_/D _14529_/Y vssd1 vssd1 vccd1 vccd1 _15467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12679_ _12679_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__xor2_1
XANTENNA__14246__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater728_A _15680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14418_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14418_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15398_ _15433_/CLK _15398_/D _14456_/Y vssd1 vssd1 vccd1 vccd1 _15398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14349_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14349_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09059__B _15364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13523__B1 _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ _08910_/A vssd1 vssd1 vccd1 vccd1 _15212_/D sky130_fd_sc_hd__clkbuf_1
X_09890_ _09889_/A _09889_/C _09977_/A vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__a21oi_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__A _15495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08841_/A _08841_/B vssd1 vssd1 vccd1 vccd1 _13914_/A sky130_fd_sc_hd__nand2_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07753__A1 _07753_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ _13880_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _15072_/D sky130_fd_sc_hd__xor2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07723_ _07723_/A vssd1 vssd1 vccd1 vccd1 _15405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1031 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ _07654_/A vssd1 vssd1 vccd1 vccd1 _15439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08419__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ _15472_/Q _07585_/A1 _07591_/S vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _15407_/Q _15391_/Q _09323_/B vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__a21o_2
XFILLER_43_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ _09254_/A _09254_/C _09254_/B vssd1 vssd1 vccd1 vccd1 _09258_/C sky130_fd_sc_hd__a21o_1
XFILLER_194_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14156__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _08292_/B _08206_/B vssd1 vssd1 vccd1 vccd1 _08231_/B sky130_fd_sc_hd__xnor2_2
XFILLER_193_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07469__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ _15571_/Q _15551_/Q vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__or2b_1
XANTENNA__08154__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08137_ _11617_/A vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__inv_2
XANTENNA__13995__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08068_ _08068_/A _11432_/B vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__xnor2_4
XFILLER_161_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1068 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _10391_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _14974_/D sky130_fd_sc_hd__xnor2_2
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput203 x_r_4[2] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13299__A_N _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 x_r_5[12] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__clkbuf_2
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__A1 _07744_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput225 x_r_5[8] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__clkbuf_1
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 x_r_6[3] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__clkbuf_2
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput247 x_r_7[13] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput258 x_r_7[9] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__clkbuf_1
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14976__D _14976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _12126_/A _11981_/B vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__nand2_2
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _14978_/Q _13836_/B vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10932_ _10931_/A _10931_/B _11127_/A vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__a21o_1
XANTENNA_input211_A x_r_5[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09432__B _15515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13651_ _13651_/A _13651_/B vssd1 vssd1 vccd1 vccd1 _13652_/B sky130_fd_sc_hd__nor2_2
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10863_ _14921_/Q _10860_/Y _10867_/B vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ _14948_/Q _12602_/B vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__and2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13582_ _13478_/A _13581_/B _13478_/B vssd1 vssd1 vccd1 vccd1 _13583_/B sky130_fd_sc_hd__a21bo_1
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _11296_/A sky130_fd_sc_hd__nor2_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15763_/CLK _15321_/D _14374_/Y vssd1 vssd1 vccd1 vccd1 _15321_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ _12533_/A _12533_/B vssd1 vssd1 vccd1 vccd1 _15613_/D sky130_fd_sc_hd__xnor2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14066__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _15268_/CLK _15252_/D _14302_/Y vssd1 vssd1 vccd1 vccd1 _15252_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12464_ _12464_/A _12464_/B vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1170 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14203_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14203_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11415_ _11414_/B _11414_/C _11414_/A vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__o21a_1
XFILLER_184_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15183_ _15775_/CLK _15183_/D _14228_/Y vssd1 vssd1 vccd1 vccd1 _15183_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08224__A2 _08223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _12395_/A _12401_/B _12401_/C vssd1 vssd1 vccd1 vccd1 _12395_/Y sky130_fd_sc_hd__nand3_1
XFILLER_153_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__inv_2
X_11346_ _11346_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__xor2_2
XFILLER_4_663 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14065_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14065_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12314__A _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _11277_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11277_/Y sky130_fd_sc_hd__nor2_1
X_13016_ _13016_/A _13016_/B _13017_/A vssd1 vssd1 vccd1 vccd1 _13016_/X sky130_fd_sc_hd__and3_1
X_10228_ _15076_/Q _15241_/Q vssd1 vssd1 vccd1 vccd1 _10230_/A sky130_fd_sc_hd__or2_1
XANTENNA_output430_A output430/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12033__B _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_475 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output528_A _15632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15047__D _15047_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__nor2_2
XFILLER_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07842__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater580_A repeater581/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ _15428_/CLK _14967_/D _14000_/Y vssd1 vssd1 vccd1 vccd1 _14967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater678_A _14526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ _14889_/A vssd1 vssd1 vccd1 vccd1 _13937_/A sky130_fd_sc_hd__buf_12
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14898_ _15729_/CLK _14898_/D _13927_/Y vssd1 vssd1 vccd1 vccd1 _14898_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _14981_/Q _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13849_/X sky130_fd_sc_hd__and3_1
XFILLER_211_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13799__B _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15519_ _15528_/CLK _15519_/D _14584_/Y vssd1 vssd1 vccd1 vccd1 _15519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09040_ _09038_/X _09045_/B vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__and2b_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_759 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14704__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_984 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09942_ _09942_/A vssd1 vssd1 vccd1 vccd1 _14965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09873_ _15187_/Q _15220_/Q vssd1 vssd1 vccd1 vccd1 _09874_/B sky130_fd_sc_hd__nand2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07726__A1 _07726_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08824_ _08824_/A _08832_/A vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__nand2_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11782__B _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08755_ _13641_/A vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__inv_2
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07706_ _15413_/Q _07706_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07707_/A sky130_fd_sc_hd__mux2_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08686_ _13491_/S _12672_/B vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08149__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07637_/A vssd1 vssd1 vccd1 vccd1 _15447_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07568_ _07568_/A vssd1 vssd1 vccd1 vccd1 _15481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09307_ _09371_/A _09307_/B vssd1 vssd1 vccd1 vccd1 _15126_/D sky130_fd_sc_hd__xor2_1
XFILLER_107_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07499_ _07499_/A vssd1 vssd1 vccd1 vccd1 _15515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09238_ _09236_/A _09236_/B _09237_/X vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__a21o_1
XFILLER_182_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _09645_/A _09169_/B vssd1 vssd1 vccd1 vccd1 _15290_/D sky130_fd_sc_hd__xnor2_1
XFILLER_135_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14614__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11200_ _11372_/A _11200_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand2_4
X_12180_ _12181_/A _12181_/B _12181_/C vssd1 vssd1 vccd1 vccd1 _12180_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__A _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11761__A2 _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__xor2_1
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input161_A x_r_1[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09427__B _15514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__A _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11062_ _14931_/Q _14997_/Q vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__or2b_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10013_ _10014_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__nor2_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14821_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input22_A x_i_1[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11692__B _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14752_/Y sky130_fd_sc_hd__inv_2
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12308_/S _12178_/A _11963_/B _11963_/C vssd1 vssd1 vccd1 vccd1 _11965_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13703_/A _13703_/B vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__xnor2_2
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _11124_/A _10915_/B vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__nand2_4
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14683_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14683_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ _11799_/A _11799_/B _11811_/B _11815_/A vssd1 vssd1 vccd1 vccd1 _11896_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13634_ _13634_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__nand2_1
XFILLER_189_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10846_ _15311_/Q vssd1 vssd1 vccd1 vccd1 _10846_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13565_ _13565_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _15603_/D sky130_fd_sc_hd__xnor2_1
X_10777_ _15787_/Q _15721_/Q vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__and2b_1
XFILLER_201_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15304_ _15592_/CLK _15304_/D _14356_/Y vssd1 vssd1 vccd1 vccd1 _15304_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11213__A _15753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12516_ _12516_/A _12516_/B _12618_/A vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__and3_1
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ _15772_/Q _13513_/A vssd1 vssd1 vccd1 vccd1 _13497_/B sky130_fd_sc_hd__or2_1
XANTENNA_output380_A output380/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output478_A _11272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15235_ _15477_/CLK _15235_/D _14284_/Y vssd1 vssd1 vccd1 vccd1 _15235_/Q sky130_fd_sc_hd__dfrtp_1
X_12447_ _12479_/A _12478_/A _12599_/A vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__or3_1
XFILLER_8_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14524__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput507 output507/A vssd1 vssd1 vccd1 vccd1 y_r_6[2] sky130_fd_sc_hd__buf_2
XFILLER_201_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput518 _15638_/Q vssd1 vssd1 vccd1 vccd1 y_r_7[12] sky130_fd_sc_hd__buf_2
X_15166_ _15775_/CLK _15166_/D _14210_/Y vssd1 vssd1 vccd1 vccd1 _15166_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12378_ _11719_/B _12378_/B vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__and2b_1
XFILLER_125_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08522__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput529 output529/A vssd1 vssd1 vccd1 vccd1 y_r_7[7] sky130_fd_sc_hd__buf_2
XFILLER_181_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14117_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11329_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__nor2_1
X_15097_ _15375_/CLK _15097_/D _14137_/Y vssd1 vssd1 vccd1 vccd1 _15097_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14048_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14048_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07708__A1 _07708_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater795_A _15594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater962_A input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08540_ _08540_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__xor2_2
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _14905_/Q vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__buf_4
XFILLER_165_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07892__A0 _15321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ _15552_/Q _07422_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15240__D _15240_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _15373_/Q _15357_/Q vssd1 vssd1 vccd1 vccd1 _09023_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14434__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09925_ _15193_/Q _09924_/Y _09920_/B vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__a21o_1
XFILLER_172_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09856_ _15064_/Q _09855_/Y _09854_/B vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08807_ _15342_/Q _15326_/Q vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__or2b_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09787_ _09562_/Y _09786_/B _09564_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__o21ai_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08738_ _08733_/X _08736_/X _08737_/X vssd1 vssd1 vccd1 vccd1 _08738_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08669_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08669_/X sky130_fd_sc_hd__or2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14609__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10700_ _10698_/X _10706_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__and2b_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11680_ _11680_/A _11680_/B _11680_/C vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__and3_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08607__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10631_ _10966_/A _10631_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12129__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13350_ _13350_/A _13356_/A _13350_/C vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__or3_1
XFILLER_195_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ _15263_/Q _15296_/Q vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__or2b_1
XFILLER_182_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12302_/A _12301_/B vssd1 vssd1 vccd1 vccd1 _15590_/D sky130_fd_sc_hd__xnor2_1
X_13281_ _13737_/B _13295_/B vssd1 vssd1 vccd1 vccd1 _13723_/B sky130_fd_sc_hd__xor2_4
XFILLER_155_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _15253_/Q _15286_/Q vssd1 vssd1 vccd1 vccd1 _10493_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14344__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07657__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15020_ _15439_/CLK _15020_/D _14056_/Y vssd1 vssd1 vccd1 vccd1 _15020_/Q sky130_fd_sc_hd__dfrtp_1
X_12232_ _12229_/Y _12230_/X _12231_/Y _12164_/A vssd1 vssd1 vccd1 vccd1 _12234_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12931__A1 _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12163_ _12238_/A _12178_/A _12308_/S vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _10886_/A _11113_/B _10886_/B vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__a21boi_2
XFILLER_122_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12094_ _12428_/A _12223_/A _12455_/C vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__or3_1
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11045_ _11039_/A _11041_/B _11039_/B vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__a21boi_1
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_754 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07392__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14804_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14804_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1018 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _15784_/CLK _15784_/D _14864_/Y vssd1 vssd1 vccd1 vccd1 _15784_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12996_ _13422_/A _13357_/B _12995_/C vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__a21oi_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14735_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14735_/Y sky130_fd_sc_hd__inv_2
X_11947_ _11947_/A _12022_/A vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__and2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14519__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07874__A0 _15330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14666_/Y sky130_fd_sc_hd__inv_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _11878_/A _11878_/B vssd1 vssd1 vccd1 vccd1 _11890_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08517__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13617_ _15375_/Q _15359_/Q vssd1 vssd1 vccd1 vccd1 _13618_/C sky130_fd_sc_hd__and2_1
X_10829_ _15307_/Q _15142_/Q vssd1 vssd1 vccd1 vccd1 _10829_/X sky130_fd_sc_hd__and2b_1
XFILLER_32_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14597_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07626__A0 _15452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13548_ _15763_/Q vssd1 vssd1 vccd1 vccd1 _13549_/A sky130_fd_sc_hd__inv_2
XFILLER_185_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater710_A _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__A _10782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ _13480_/C _13480_/B _13581_/A vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__a21boi_1
XANTENNA_repeater808_A _15581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14254__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ _15727_/CLK _15218_/D _14266_/Y vssd1 vssd1 vccd1 vccd1 _15218_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__07567__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput304 output304/A vssd1 vssd1 vccd1 vccd1 y_i_2[3] sky130_fd_sc_hd__buf_2
XANTENNA__08252__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput315 _15673_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[13] sky130_fd_sc_hd__buf_2
Xoutput326 _15668_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[8] sky130_fd_sc_hd__buf_2
XFILLER_154_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput337 _11305_/Y vssd1 vssd1 vccd1 vccd1 y_i_4[2] sky130_fd_sc_hd__buf_2
X_15149_ _15394_/CLK _15149_/D _14192_/Y vssd1 vssd1 vccd1 vccd1 _15149_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput348 _15688_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[12] sky130_fd_sc_hd__buf_2
Xoutput359 _15683_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[7] sky130_fd_sc_hd__buf_2
XFILLER_82_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07971_ _10722_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _07971_/Y sky130_fd_sc_hd__nor2_2
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09710_ _15059_/Q _15092_/Q vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09083__A _15497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ _09639_/A _09639_/B _09640_/X vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15813__A _15813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _15437_/Q _15421_/Q vssd1 vssd1 vccd1 vccd1 _09572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08523_ _08603_/B _08538_/B _12688_/A vssd1 vssd1 vccd1 vccd1 _08524_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_971 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14429__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11661__A1 _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _08728_/B _12945_/A vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07405_ _07405_/A vssd1 vssd1 vccd1 vccd1 _15565_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _12654_/A vssd1 vssd1 vccd1 vccd1 _08385_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12891__B _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__A2 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14164__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ _15370_/Q _15354_/Q vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07477__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09908_ _15192_/Q _15225_/Q vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12412__A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09839_ _15093_/Q _15060_/Q vssd1 vssd1 vccd1 vccd1 _09840_/C sky130_fd_sc_hd__or2b_1
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12131__B _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12850_ _15762_/Q vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__inv_2
XFILLER_98_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input124_A x_i_7[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _12308_/S _12178_/A vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__or2_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12781_/A _12781_/B vssd1 vssd1 vccd1 vccd1 _12781_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14339__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_695 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13243__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14520_/Y sky130_fd_sc_hd__inv_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14451_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _12122_/A _11977_/A _11663_/C vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__and3_1
XFILLER_35_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ _15769_/Q _13576_/B vssd1 vssd1 vccd1 vccd1 _13574_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07608__A0 _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ _10614_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _14998_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14382_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14382_/Y sky130_fd_sc_hd__inv_2
X_11594_ _11797_/A _08009_/C _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11594_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_161_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09073__A2 _15478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11698__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13333_ _13333_/A _13333_/B _13333_/C vssd1 vssd1 vccd1 vccd1 _13335_/A sky130_fd_sc_hd__or3_1
X_10545_ _10545_/A _10551_/A vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__and2_1
XANTENNA__14074__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_130_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15508_/CLK sky130_fd_sc_hd__clkbuf_16
X_13264_ _13264_/A _13308_/A vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__nor2_1
X_10476_ _15163_/Q vssd1 vssd1 vccd1 vccd1 _10476_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ _15509_/CLK _15003_/D _14037_/Y vssd1 vssd1 vccd1 vccd1 _15003_/Q sky130_fd_sc_hd__dfrtp_1
X_12215_ _12466_/A _12216_/B vssd1 vssd1 vccd1 vccd1 _12215_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13195_ _13195_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13196_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13502__A_N _13790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12146_ _12088_/A _12088_/B _12087_/A vssd1 vssd1 vccd1 vccd1 _12209_/B sky130_fd_sc_hd__a21oi_1
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output343_A output343/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _12186_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__and2_1
Xrepeater807 _15582_/Q vssd1 vssd1 vccd1 vccd1 output425/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08336__A1 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater818 input99/X vssd1 vssd1 vccd1 vccd1 _07543_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08336__B2 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater829 repeater830/X vssd1 vssd1 vccd1 vccd1 _07453_/A1 sky130_fd_sc_hd__buf_4
X_11028_ _14924_/Q _14990_/Q vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output510_A output510/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07850__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__B _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _13681_/B _12979_/B vssd1 vssd1 vccd1 vccd1 _13549_/B sky130_fd_sc_hd__xnor2_4
X_15767_ _15774_/CLK _15767_/D _14846_/Y vssd1 vssd1 vccd1 vccd1 _15767_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater758_A _15643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14249__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14718_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14718_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08247__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15698_ _15770_/CLK _15698_/D _14773_/Y vssd1 vssd1 vccd1 vccd1 _15698_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14649_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14649_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_838 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08170_ _12312_/S _11471_/B vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__xnor2_1
XFILLER_177_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15460_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09078__A _15496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14712__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ _14921_/Q _15775_/Q vssd1 vssd1 vccd1 vccd1 _11105_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07885_ _07885_/A vssd1 vssd1 vccd1 vccd1 _15325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09624_ _15444_/Q _15428_/Q vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__and2b_1
XFILLER_46_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09555_ _15432_/Q _15416_/Q vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14159__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08506_/X sky130_fd_sc_hd__or2_1
XANTENNA__07838__A0 _15348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _09486_/A _09486_/B vssd1 vssd1 vccd1 vccd1 _15281_/D sky130_fd_sc_hd__nor2_2
XFILLER_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13998__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _08437_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _08459_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07996__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _15046_/Q vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08299_ _11658_/A _11687_/A _11617_/A _11584_/A _08298_/X vssd1 vssd1 vccd1 vccd1
+ _08299_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_112_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ _10324_/A _10326_/B _10324_/B vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__a21boi_2
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10261_ _10260_/A _10260_/B _11414_/A vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__a21o_1
XFILLER_127_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14622__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12000_ _12079_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__or2_1
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _09688_/Y _15218_/Q _11392_/B vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14979__D _14979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input241_A x_r_6[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12902_ _12902_/A _12902_/B _12900_/Y vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__or3b_1
X_13882_ _15336_/Q _15320_/Q _13881_/X vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__a21oi_2
XFILLER_47_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15621_ _15724_/CLK _15621_/D _14692_/Y vssd1 vssd1 vccd1 vccd1 _15621_/Q sky130_fd_sc_hd__dfrtp_1
X_12833_ _12906_/A _12833_/B vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__and2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14069__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _13056_/C _12764_/B vssd1 vssd1 vccd1 vccd1 _12775_/A sky130_fd_sc_hd__xnor2_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15571_/CLK _15552_/D _14618_/Y vssd1 vssd1 vccd1 vccd1 _15552_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ _11728_/A _12390_/A vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__or2_1
X_14503_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14503_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15483_/CLK _15483_/D _14546_/Y vssd1 vssd1 vccd1 vccd1 _15483_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _13645_/A _13645_/B vssd1 vssd1 vccd1 vccd1 _13649_/B sky130_fd_sc_hd__xnor2_4
XFILLER_70_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11646_ _11646_/A _11646_/B vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__xnor2_2
X_14434_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output293_A output293/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 x_i_0[5] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput25 x_i_1[15] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14365_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14365_/Y sky130_fd_sc_hd__inv_2
Xinput36 x_i_2[10] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
X_11577_ _11577_/A vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_103_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15341_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 x_i_2[6] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 x_i_3[1] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
X_13316_ _13277_/X _13316_/B _13316_/C vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__and3b_1
XANTENNA__11221__A _15032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 x_i_4[11] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_4
XFILLER_143_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10528_ _15290_/Q _15257_/Q vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__and2b_1
XFILLER_196_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output460_A _15600_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14296_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14296_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13247_ _13247_/A _13247_/B vssd1 vssd1 vccd1 vccd1 _13248_/B sky130_fd_sc_hd__nand2_1
X_10459_ _10459_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14532__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09626__A _15541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ _13352_/A _15052_/Q vssd1 vssd1 vccd1 vccd1 _13250_/B sky130_fd_sc_hd__and2_1
XANTENNA__08530__A _08530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12129_ _12247_/A _12244_/A vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13148__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater604 repeater605/X vssd1 vssd1 vccd1 vccd1 output410/A sky130_fd_sc_hd__buf_4
Xrepeater615 _11361_/Y vssd1 vssd1 vccd1 vccd1 output442/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater626 _10738_/Y vssd1 vssd1 vccd1 vccd1 output407/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater637 _11026_/Y vssd1 vssd1 vccd1 vccd1 output269/A sky130_fd_sc_hd__clkbuf_2
Xrepeater648 _07975_/X vssd1 vssd1 vccd1 vccd1 _15810_/A sky130_fd_sc_hd__buf_2
XANTENNA_repeater875_A input253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater659 _14787_/A vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__buf_4
X_07670_ _07670_/A vssd1 vssd1 vccd1 vccd1 _15431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09340_ _09340_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _15133_/D sky130_fd_sc_hd__xor2_4
XFILLER_179_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _15249_/D sky130_fd_sc_hd__xnor2_1
XFILLER_205_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14707__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ _12008_/A vssd1 vssd1 vccd1 vccd1 _11842_/C sky130_fd_sc_hd__inv_2
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08192_/A sky130_fd_sc_hd__xor2_1
XFILLER_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _08071_/Y _08083_/A _08081_/X _08094_/B _08094_/A vssd1 vssd1 vccd1 vccd1
+ _08086_/B sky130_fd_sc_hd__a32o_1
XFILLER_88_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13698__A_N _13827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14442__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07755__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _08986_/A _08986_/B _13594_/A vssd1 vssd1 vccd1 vccd1 _08988_/A sky130_fd_sc_hd__nor3_1
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07937_ _15086_/Q vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__inv_2
XFILLER_180_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07868_ _15333_/Q input195/X _07900_/S vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A vssd1 vssd1 vccd1 vccd1 _15180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07799_ _15367_/Q _07799_/A1 _07803_/S vssd1 vssd1 vccd1 vccd1 _07800_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ _15430_/Q _15414_/Q vssd1 vssd1 vccd1 vccd1 _09545_/A sky130_fd_sc_hd__and2b_1
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13224__C _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09469_ _09469_/A vssd1 vssd1 vccd1 vccd1 _15278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14617__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _11498_/Y _08316_/A _08316_/B _11499_/Y vssd1 vssd1 vccd1 vccd1 _11501_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_169_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12480_ _12464_/B _12479_/Y _12604_/A _12601_/A vssd1 vssd1 vccd1 vccd1 _12488_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__A1 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input191_A x_r_3[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14150_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_898 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11362_ _11172_/A _11361_/B _11172_/B vssd1 vssd1 vccd1 vccd1 _11363_/B sky130_fd_sc_hd__a21boi_4
XFILLER_165_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A _13044_/B vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__or2b_1
XFILLER_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11976__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10313_ _15124_/Q _15157_/Q vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__nand2_1
X_14081_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__inv_2
X_11293_ _11292_/A _11292_/B _10778_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14352__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ _13109_/B _12784_/C _13220_/A vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11695__B _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A x_i_3[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _11411_/A _10244_/B vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__nand2_2
XFILLER_191_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08350__A _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10852_/A sky130_fd_sc_hd__nor2_2
XFILLER_26_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14983_ _15773_/CLK _14983_/D _14016_/Y vssd1 vssd1 vccd1 vccd1 _14983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11915__S _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13934_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13415__B _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ _13865_/A _13868_/B vssd1 vssd1 vccd1 vccd1 _15674_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output306_A output306/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13599__A1 _15368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ _15774_/CLK _15604_/D _14674_/Y vssd1 vssd1 vccd1 vccd1 _15604_/Q sky130_fd_sc_hd__dfrtp_1
X_12816_ _13357_/B _13201_/A vssd1 vssd1 vccd1 vccd1 _12893_/C sky130_fd_sc_hd__xor2_2
XFILLER_76_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13796_ _13789_/A _13863_/A _13788_/A vssd1 vssd1 vccd1 vccd1 _13797_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ _15563_/CLK _15535_/D _14600_/Y vssd1 vssd1 vccd1 vccd1 _15535_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _14920_/Q _12791_/B vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__A_N _15476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14527__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12750_/A _12750_/B vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__xor2_1
X_15466_ _15558_/CLK _15466_/D _14528_/Y vssd1 vssd1 vccd1 vccd1 _15466_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11629_ _12144_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _11697_/C sky130_fd_sc_hd__xor2_2
X_14417_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14417_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater623_A _11359_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ _15399_/CLK _15397_/D _14455_/Y vssd1 vssd1 vccd1 vccd1 _15397_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_204_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14348_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10790__A _10790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14262__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13523__A1 _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__S _07575_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _15348_/Q _15332_/Q vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__or2_1
XFILLER_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08770_/Y _15319_/Q _08768_/B vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__a21o_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07722_ _15405_/Q _07722_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07653_ _15439_/Q _07653_/A1 _07687_/S vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09972__A1_N _15186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1043 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07584_ _07584_/A vssd1 vssd1 vccd1 vccd1 _15473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _15129_/D sky130_fd_sc_hd__nor2_1
XFILLER_40_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14437__A _14439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09254_ _09254_/A _09254_/B _09254_/C vssd1 vssd1 vccd1 vccd1 _09254_/X sky130_fd_sc_hd__and3_1
XFILLER_22_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08205_ _11467_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08206_/B sky130_fd_sc_hd__nand2_1
XFILLER_194_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09185_ _15551_/Q _15571_/Q vssd1 vssd1 vccd1 vccd1 _09187_/A sky130_fd_sc_hd__or2b_1
XFILLER_147_640 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08136_ _11467_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07441__A1 _07441_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08290_/B _08118_/B _08066_/Y vssd1 vssd1 vccd1 vccd1 _11432_/B sky130_fd_sc_hd__a21o_2
XFILLER_175_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14172__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07485__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08170__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_955 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 x_r_4[3] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__clkbuf_1
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 x_r_5[13] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput226 x_r_5[9] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__08941__A1 _15463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 x_r_6[4] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_4
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 x_r_7[14] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08969_ _08967_/A _08967_/B _08968_/X vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__a21o_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11980_ _11980_/A _11980_/B _11978_/Y vssd1 vssd1 vccd1 vccd1 _11981_/B sky130_fd_sc_hd__or3b_1
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09497__A2 _15509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_671 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _10931_/A _10931_/B _11127_/A vssd1 vssd1 vccd1 vccd1 _10931_/X sky130_fd_sc_hd__and3_1
XFILLER_205_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input204_A x_r_4[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862_ _10861_/Y _15775_/Q _11105_/B vssd1 vssd1 vccd1 vccd1 _10867_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13650_ _13649_/A _13649_/B _13638_/B _13638_/A vssd1 vssd1 vccd1 vccd1 _13651_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _15686_/D sky130_fd_sc_hd__xor2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _15607_/D sky130_fd_sc_hd__xnor2_1
X_10793_ _15789_/Q _15723_/Q vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__and2b_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14347__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13251__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12532_ _12530_/X _12529_/B _12531_/X vssd1 vssd1 vccd1 vccd1 _12533_/B sky130_fd_sc_hd__a21o_1
X_15320_ _15352_/CLK _15320_/D _14373_/Y vssd1 vssd1 vccd1 vccd1 _15320_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _14947_/Q _12463_/B _12463_/C vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__nand3_1
X_15251_ _15268_/CLK _15251_/D _14301_/Y vssd1 vssd1 vccd1 vccd1 _15251_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14202_/Y sky130_fd_sc_hd__inv_2
X_11414_ _11414_/A _11414_/B _11414_/C vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__nor3_1
X_15182_ _15775_/CLK _15182_/D _14227_/Y vssd1 vssd1 vccd1 vccd1 _15182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_1182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12394_ _12401_/B _12401_/C _12395_/A vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__a21oi_1
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14133_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14133_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07432__A1 _07432_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _11344_/A _11344_/B _11076_/B vssd1 vssd1 vccd1 vccd1 _11346_/B sky130_fd_sc_hd__a21o_1
XFILLER_181_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14082__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_675 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14064_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14064_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11276_ _11275_/B _11275_/C _11275_/A vssd1 vssd1 vccd1 vccd1 _11277_/B sky130_fd_sc_hd__a21oi_1
XFILLER_180_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _13015_/A _13069_/B vssd1 vssd1 vccd1 vccd1 _13023_/A sky130_fd_sc_hd__xor2_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _15764_/D sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_88_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14810__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__C _13713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__C _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10158_ _15312_/Q _15147_/Q vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__and2b_1
XANTENNA_output423_A _15580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_131_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14966_ _15727_/CLK _14966_/D _13999_/Y vssd1 vssd1 vccd1 vccd1 _14966_/Q sky130_fd_sc_hd__dfrtp_1
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _14984_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14889_/A sky130_fd_sc_hd__buf_12
XFILLER_78_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12492__A1 _12262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14897_ _15729_/CLK _14897_/D _13926_/Y vssd1 vssd1 vccd1 vccd1 _14897_/Q sky130_fd_sc_hd__dfrtp_1
X_13848_ _13848_/A _13848_/B vssd1 vssd1 vccd1 vccd1 _15671_/D sky130_fd_sc_hd__xor2_1
XFILLER_74_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_26_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater838_A input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ _13775_/A _13862_/B _13778_/X vssd1 vssd1 vccd1 vccd1 _13779_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__14257__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15518_ _15563_/CLK _15518_/D _14583_/Y vssd1 vssd1 vccd1 vccd1 _15518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_15449_ _15493_/CLK _15449_/D _14510_/Y vssd1 vssd1 vccd1 vccd1 _15449_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15118__RESET_B _14160_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _09939_/X _09946_/B vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__and2b_1
XFILLER_132_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15238__D _15238_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15816__A _15816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _15187_/Q _15220_/Q vssd1 vssd1 vccd1 vccd1 _09872_/Y sky130_fd_sc_hd__nor2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14720__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _15345_/Q _15329_/Q vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__or2b_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13336__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08754_ _14938_/Q _13808_/A vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07705_ _07705_/A vssd1 vssd1 vccd1 vccd1 _15414_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08685_/A _12667_/C vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__xnor2_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08149__B _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _15447_/Q input11/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07567_ _15481_/Q input45/X _07579_/S vssd1 vssd1 vccd1 vccd1 _07568_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14167__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09306_ _15403_/Q _15387_/Q _09305_/X vssd1 vssd1 vccd1 vccd1 _09307_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07498_ _15515_/Q input31/X _07536_/S vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ _15499_/Q _15483_/Q vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__and2b_1
XFILLER_186_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ _09161_/Y _09166_/B _09163_/B vssd1 vssd1 vccd1 vccd1 _09169_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08119_ _08323_/A _08323_/B _08271_/A vssd1 vssd1 vccd1 vccd1 _08119_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07414__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09099_ _15499_/Q _15483_/Q _09098_/X vssd1 vssd1 vccd1 vccd1 _09100_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08612__B _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _14965_/Q _14899_/Q _11129_/B vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__a21o_1
XFILLER_135_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11333_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/Y sky130_fd_sc_hd__xnor2_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input154_A x_r_1[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14630__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _10383_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__nand2_1
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14820_/Y sky130_fd_sc_hd__inv_2
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A x_i_0[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14751_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _11882_/A _11963_/B _11963_/C vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__and3b_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15741_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13702_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__or2b_1
X_10914_ _14963_/Q _14897_/Q vssd1 vssd1 vccd1 vccd1 _10915_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _11894_/A _11894_/B vssd1 vssd1 vccd1 vccd1 _11953_/B sky130_fd_sc_hd__xor2_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14701_/A sky130_fd_sc_hd__buf_12
XFILLER_205_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10845_ _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _14915_/D sky130_fd_sc_hd__nor2_1
X_13633_ _14971_/Q vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__inv_2
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15611__D _15611_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14077__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10776_ _15721_/Q _15787_/Q vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__and2b_1
XFILLER_13_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__D1 _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _13564_/A _13564_/B vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15303_ _15592_/CLK _15303_/D _14355_/Y vssd1 vssd1 vccd1 vccd1 _15303_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07653__A1 _07653_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ _12516_/A _12516_/B _12618_/A vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__a21oi_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13495_ _15772_/Q _13513_/A vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__nand2_1
XFILLER_200_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14805__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12446_ _12479_/A _12478_/A _12599_/A vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__o21ai_1
X_15234_ _15493_/CLK _15234_/D _14283_/Y vssd1 vssd1 vccd1 vccd1 _15234_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output373_A output373/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput508 output508/A vssd1 vssd1 vccd1 vccd1 y_r_6[3] sky130_fd_sc_hd__buf_2
X_12377_ _12375_/A _12582_/A _12376_/X vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__a21o_1
XFILLER_172_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15165_ _15180_/CLK _15165_/D _14209_/Y vssd1 vssd1 vccd1 vccd1 _15165_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput519 output519/A vssd1 vssd1 vccd1 vccd1 y_r_7[13] sky130_fd_sc_hd__buf_2
XANTENNA__08522__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14116_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14116_/Y sky130_fd_sc_hd__inv_2
X_11328_ _11327_/B _11327_/C _11327_/A vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__a21oi_1
XFILLER_10_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15096_ _15375_/CLK _15096_/D _14136_/Y vssd1 vssd1 vccd1 vccd1 _15096_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14047_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14047_/Y sky130_fd_sc_hd__inv_2
X_11259_ _11259_/A _11259_/B _11259_/C vssd1 vssd1 vccd1 vccd1 _11261_/A sky130_fd_sc_hd__and3_1
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14540__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09634__A _15563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__B _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12783__A_N _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater690_A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater788_A _15604_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _15790_/CLK _14949_/D _13981_/Y vssd1 vssd1 vccd1 vccd1 _14949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater955_A input141/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12995__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ _14907_/Q vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__buf_6
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _07421_/A vssd1 vssd1 vccd1 vccd1 _15553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07892__A1 _07892_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07644__A1 _07644_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14715__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ _09022_/A vssd1 vssd1 vccd1 vccd1 _13612_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09924_ _15226_/Q vssd1 vssd1 vccd1 vccd1 _09924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14450__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11793__B _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__A _15431_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _15097_/Q vssd1 vssd1 vccd1 vccd1 _09855_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input7_A x_i_0[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ _13895_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _15158_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08737_ _08734_/Y _08735_/X _08722_/Y _08723_/X vssd1 vssd1 vccd1 vccd1 _08737_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15699_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_855 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08668_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _08671_/A sky130_fd_sc_hd__xnor2_4
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_814 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _07619_/A vssd1 vssd1 vccd1 vccd1 _15456_/D sky130_fd_sc_hd__clkbuf_1
X_08599_ _08599_/A _08619_/A vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__nand2_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10630_ _15268_/Q _15169_/Q vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__or2b_1
XFILLER_197_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12129__B _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10561_ _10561_/A vssd1 vssd1 vccd1 vccd1 _15031_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14625__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _12299_/Y _12564_/B _12270_/B vssd1 vssd1 vccd1 vccd1 _12301_/B sky130_fd_sc_hd__o21ai_2
XFILLER_10_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09719__A _15061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ _13280_/A _13280_/B vssd1 vssd1 vccd1 vccd1 _13295_/B sky130_fd_sc_hd__xnor2_4
XFILLER_155_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _15251_/Q _10490_/Y _10496_/B vssd1 vssd1 vccd1 vccd1 _15021_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12231_ _12231_/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09438__B _15515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12162_ _12308_/S _12238_/A vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12931__A2 _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11113_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12093_ _12451_/B _12105_/B vssd1 vssd1 vccd1 vccd1 _12455_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__14360__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11044_ _11042_/Y _11044_/B vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__and2b_1
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_766 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _15790_/CLK _15783_/D _14863_/Y vssd1 vssd1 vccd1 vccd1 _15783_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15727_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12995_ _13422_/A _13357_/B _12995_/C vssd1 vssd1 vccd1 vccd1 _13192_/B sky130_fd_sc_hd__and3_1
XFILLER_80_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14741_/A vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11946_ _11945_/A _11945_/B _12547_/A vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__o21ai_2
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07874__A1 input135/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13431__A_N _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14665_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14665_/Y sky130_fd_sc_hd__inv_2
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11877_ _11877_/A vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__inv_2
XFILLER_162_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _13616_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _15096_/D sky130_fd_sc_hd__nor2_1
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ _10828_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _14911_/D sky130_fd_sc_hd__xor2_2
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output490_A _15612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1090 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07626__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13547_ _13547_/A _13547_/B vssd1 vssd1 vccd1 vccd1 _15599_/D sky130_fd_sc_hd__xor2_2
X_10759_ _15718_/Q _15784_/Q vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__or2_1
XANTENNA__14535__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07848__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13478_ _13478_/A _13478_/B vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08533__A _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15217_ _15460_/CLK _15217_/D _14265_/Y vssd1 vssd1 vccd1 vccd1 _15217_/Q sky130_fd_sc_hd__dfrtp_1
X_12429_ _12430_/B _12430_/C _12455_/B vssd1 vssd1 vccd1 vccd1 _12440_/C sky130_fd_sc_hd__o21a_1
XANTENNA_repeater703_A _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput305 output305/A vssd1 vssd1 vccd1 vccd1 y_i_2[4] sky130_fd_sc_hd__buf_2
XANTENNA__12055__A _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__B _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput316 _15674_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[14] sky130_fd_sc_hd__buf_2
XFILLER_99_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput327 _15669_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[9] sky130_fd_sc_hd__buf_2
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput338 _11308_/X vssd1 vssd1 vccd1 vccd1 y_i_4[3] sky130_fd_sc_hd__buf_2
X_15148_ _15394_/CLK _15148_/D _14191_/Y vssd1 vssd1 vccd1 vccd1 _15148_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput349 _15689_/Q vssd1 vssd1 vccd1 vccd1 y_i_5[13] sky130_fd_sc_hd__buf_2
XFILLER_114_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _15775_/Q _15709_/Q vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ _15081_/CLK _15079_/D _14118_/Y vssd1 vssd1 vccd1 vccd1 _15079_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14270__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1072 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09640_ _15565_/Q _15545_/Q vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__and2b_1
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09571_ _09788_/A _09571_/B vssd1 vssd1 vccd1 vccd1 _15175_/D sky130_fd_sc_hd__xor2_1
XFILLER_27_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15439_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_208_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08522_ _12780_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__xor2_1
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08453_ _13012_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08455_/B sky130_fd_sc_hd__nor2_1
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07404_ _15565_/Q _07404_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08384_ _12881_/A _12654_/A _08384_/C vssd1 vssd1 vccd1 vccd1 _08410_/B sky130_fd_sc_hd__and3_1
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14445__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ _09003_/Y _09005_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__nand2b_1
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09790__A1 _15436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14180__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _15192_/Q _15225_/Q vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__or2_1
XFILLER_154_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09838_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07553__A0 _15488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09769_ _09767_/A _09863_/A _09768_/Y vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_38_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15808_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _12308_/S _12178_/A vssd1 vssd1 vccd1 vccd1 _11882_/A sky130_fd_sc_hd__nand2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input117_A x_i_7[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12805_/B sky130_fd_sc_hd__nand2_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11707_/A _11707_/B _11730_/X vssd1 vssd1 vccd1 vccd1 _11863_/B sky130_fd_sc_hd__a21bo_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14450_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14450_/Y sky130_fd_sc_hd__inv_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _12178_/A _12055_/A vssd1 vssd1 vccd1 vccd1 _11663_/C sky130_fd_sc_hd__xor2_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13401_ _13401_/A _13747_/B vssd1 vssd1 vccd1 vccd1 _13576_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07608__A1 input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ _10612_/B _10612_/C _10612_/A vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__o21a_1
X_11593_ _11797_/A _11876_/A vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__nor2_1
X_14381_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14381_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14355__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_552 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13332_ _13332_/A _13375_/A vssd1 vssd1 vccd1 vccd1 _13333_/C sky130_fd_sc_hd__xnor2_1
X_10544_ _10543_/A _10543_/C _10606_/A vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_input82_A x_i_4[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _14899_/D sky130_fd_sc_hd__nor2_1
X_13263_ _13263_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _13308_/A sky130_fd_sc_hd__and2_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15002_ _15509_/CLK _15002_/D _14036_/Y vssd1 vssd1 vccd1 vccd1 _15002_/Q sky130_fd_sc_hd__dfrtp_2
X_12214_ _12214_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__nor2_2
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13194_ _13195_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13270_/B sky130_fd_sc_hd__or2_1
XFILLER_159_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12145_ _12207_/B _12145_/B vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__nand2_1
XFILLER_29_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14090__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _12075_/A _12075_/B _12075_/C vssd1 vssd1 vccd1 vccd1 _12077_/B sky130_fd_sc_hd__o21ai_1
XFILLER_110_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output336_A output336/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater808 _15581_/Q vssd1 vssd1 vccd1 vccd1 output424/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater819 input98/X vssd1 vssd1 vccd1 vccd1 _07459_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__A _11219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ _14924_/Q _14990_/Q vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__or2_1
XFILLER_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output503_A _11237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15391_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12976__C _12976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15774_/CLK _15766_/D _14845_/Y vssd1 vssd1 vccd1 vccd1 _15766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ _13677_/C _12916_/B _12912_/A vssd1 vssd1 vccd1 vccd1 _12979_/B sky130_fd_sc_hd__o21ai_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14717_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14717_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13153__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11929_ _12011_/B _11929_/B vssd1 vssd1 vccd1 vccd1 _11931_/C sky130_fd_sc_hd__or2_1
X_15697_ _15774_/CLK _15697_/D _14772_/Y vssd1 vssd1 vccd1 vccd1 _15697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08247__B _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14648_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater820_A input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14579_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14579_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14265__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater918_A input190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09078__B _15480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_839 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07953_ _07953_/A vssd1 vssd1 vccd1 vccd1 _15792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15246__D _15246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07884_ _15325_/Q input145/X _07892_/S vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09623_ _09812_/A _09623_/B vssd1 vssd1 vccd1 vccd1 _15183_/D sky130_fd_sc_hd__xnor2_1
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _09552_/Y _09554_/B vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__nand2b_1
XFILLER_197_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08552_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07838__A1 input201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ _09484_/A _09484_/B _09532_/A vssd1 vssd1 vccd1 vccd1 _09486_/B sky130_fd_sc_hd__o21a_1
XFILLER_102_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08157__B _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08436_ _08441_/A _08399_/B _13201_/A vssd1 vssd1 vccd1 vccd1 _08437_/B sky130_fd_sc_hd__o21bai_1
XFILLER_178_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08367_ _13357_/B _08376_/B vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__xnor2_2
XFILLER_196_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14175__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09269__A _15507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _11584_/A _11617_/A _11491_/A _11458_/A _08297_/Y vssd1 vssd1 vccd1 vccd1
+ _08298_/X sky130_fd_sc_hd__a221o_1
XFILLER_194_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10260_ _10260_/A _10260_/B _11414_/A vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__and3_1
XFILLER_152_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10191_ _15218_/Q _11392_/B vssd1 vssd1 vccd1 vccd1 _10191_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1081 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13950_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13950_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input234_A x_r_6[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12901_ _12902_/A _12902_/B _12900_/Y vssd1 vssd1 vccd1 vccd1 _13016_/A sky130_fd_sc_hd__o21bai_1
XFILLER_115_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13881_ _15336_/Q _15320_/Q _13880_/B vssd1 vssd1 vccd1 vccd1 _13881_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _15724_/CLK _15620_/D _14691_/Y vssd1 vssd1 vccd1 vccd1 _15620_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _12832_/A _12832_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _12833_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15571_/CLK _15551_/D _14617_/Y vssd1 vssd1 vccd1 vccd1 _15551_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _13057_/A _13057_/B vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__nand2_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14502_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11714_ _11714_/A _11714_/B vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__xnor2_2
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _15500_/CLK _15482_/D _14545_/Y vssd1 vssd1 vccd1 vccd1 _15482_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _13645_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14433_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11645_ _11866_/A _11865_/C _11866_/B _11570_/A vssd1 vssd1 vccd1 vccd1 _11646_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14085__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11502__A _15727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 x_i_0[6] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
X_14364_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14364_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11576_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11577_/A sky130_fd_sc_hd__and2_1
XFILLER_167_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 x_i_1[1] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output286_A _15645_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 x_i_2[11] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 x_i_2[7] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13315_ _13315_/A _13315_/B vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__xnor2_2
Xinput59 x_i_3[2] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
X_10527_ _10527_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10602_/A sky130_fd_sc_hd__nand2_1
X_14295_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14295_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14813__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10458_ _10459_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _14895_/D sky130_fd_sc_hd__xor2_1
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13246_ _13246_/A _13245_/X vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__or2b_2
XFILLER_182_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12889__A1 _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output453_A output453/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12333__A _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ _13177_/A _13177_/B vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__nand2_1
X_10389_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ _12128_/A _12128_/B vssd1 vssd1 vccd1 vccd1 _12466_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__13148__B _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater605 _10753_/Y vssd1 vssd1 vccd1 vccd1 repeater605/X sky130_fd_sc_hd__buf_2
X_12059_ _12059_/A _12059_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__xor2_4
Xrepeater616 _11261_/Y vssd1 vssd1 vccd1 vccd1 output475/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater627 _11357_/Y vssd1 vssd1 vccd1 vccd1 output440/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater638 _10869_/Y vssd1 vssd1 vccd1 vccd1 output303/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater649 _07971_/Y vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater770_A _15628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater868_A repeater869/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15749_ _15749_/CLK _15749_/D _14827_/Y vssd1 vssd1 vccd1 vccd1 _15749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09270_ _09269_/Y _15491_/Q _09268_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08221_ _15013_/Q vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__buf_4
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08174_/B sky130_fd_sc_hd__nor2_1
XFILLER_165_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08083_ _08083_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15553_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__14723__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ _15367_/Q _15351_/Q vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _07936_/A vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07771__S _07795_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ _07867_/A vssd1 vssd1 vccd1 vccd1 _15334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _09604_/X _09611_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13074__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08168__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07798_ _07798_/A vssd1 vssd1 vccd1 vccd1 _15368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ _15413_/Q vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__inv_2
XFILLER_25_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09466_/X _09473_/B vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__and2b_1
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ _13422_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09399_ _09398_/A _09398_/C _09398_/B vssd1 vssd1 vccd1 vccd1 _09400_/B sky130_fd_sc_hd__a21oi_1
XFILLER_196_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11430_ _11430_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _15742_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__12032__A2 _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11361_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14633__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input184_A x_r_3[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _15124_/Q _15157_/Q vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__or2_1
XFILLER_138_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13100_ _13100_/A _13100_/B _13100_/C vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__nand3_2
XFILLER_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11292_ _11292_/A _11292_/B vssd1 vssd1 vccd1 vccd1 _11292_/X sky130_fd_sc_hd__xor2_2
X_14080_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14080_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _13319_/A vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__inv_2
XFILLER_69_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10243_ _15078_/Q _15243_/Q vssd1 vssd1 vccd1 vccd1 _10244_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10174_ _15314_/Q _15149_/Q vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__and2b_1
XANTENNA_input45_A x_i_2[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14982_ _15773_/CLK _14982_/D _14015_/Y vssd1 vssd1 vccd1 vccd1 _14982_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_980 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07681__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__A _09462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13933_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15614__D _15614_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13864_ _13863_/B _13863_/C _13863_/A vssd1 vssd1 vccd1 vccd1 _13868_/B sky130_fd_sc_hd__o21a_1
X_15603_ _15771_/CLK _15603_/D _14673_/Y vssd1 vssd1 vccd1 vccd1 _15603_/Q sky130_fd_sc_hd__dfrtp_2
X_12815_ _13203_/A _13273_/A vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__nand2_1
X_13795_ _14985_/Q _13871_/B vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__xor2_2
XANTENNA__14808__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _15563_/CLK _15534_/D _14599_/Y vssd1 vssd1 vccd1 vccd1 _15534_/Q sky130_fd_sc_hd__dfrtp_1
X_12746_ _12746_/A _12784_/C vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__xnor2_1
XFILLER_187_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13431__B _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15465_ _15477_/CLK _15465_/D _14527_/Y vssd1 vssd1 vccd1 vccd1 _15465_/Q sky130_fd_sc_hd__dfrtp_1
X_12677_ _13431_/B _12743_/B vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14416_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__inv_2
X_11628_ _11928_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15396_ _15575_/CLK _15396_/D _14454_/Y vssd1 vssd1 vccd1 vccd1 _15396_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14347_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14347_/Y sky130_fd_sc_hd__inv_2
X_11559_ _11559_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14543__A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07856__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14278_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14278_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13229_ _13330_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13230_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater985_A input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08770_ _15335_/Q vssd1 vssd1 vccd1 vccd1 _08770_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07721_ _07721_/A vssd1 vssd1 vccd1 vccd1 _15406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07652_ _07652_/A vssd1 vssd1 vccd1 vccd1 _15440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07583_ _15473_/Q input70/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14718__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09322_ _09321_/A _09321_/C _09382_/A vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__o21a_1
XFILLER_40_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09253_ _09253_/A vssd1 vssd1 vccd1 vccd1 _15244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12238__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08204_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08231_/A sky130_fd_sc_hd__xor2_2
X_09184_ _09654_/A _09188_/B vssd1 vssd1 vccd1 vccd1 _15293_/D sky130_fd_sc_hd__xor2_1
XFILLER_21_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13060__C _13062_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ _08223_/B vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__buf_8
XFILLER_181_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14453__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08066_ _08066_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput205 x_r_4[4] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput216 x_r_5[14] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput227 x_r_6[0] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__08941__A2 _15447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 x_r_6[5] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08968_ _08968_/A _15457_/Q vssd1 vssd1 vccd1 vccd1 _08968_/X sky130_fd_sc_hd__and2_1
Xinput249 x_r_7[15] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_1
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07919_ _07919_/A vssd1 vssd1 vccd1 vccd1 _15251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_609 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08899_ _08899_/A _08907_/A vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater980 repeater981/X vssd1 vssd1 vccd1 vccd1 _07526_/A1 sky130_fd_sc_hd__buf_4
X_10930_ _10930_/A _10938_/A vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10221__A _15075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ _14921_/Q vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14628__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ _12445_/B _12599_/B _12443_/Y vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__a21o_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13579_/A _13579_/B _15770_/Q _13451_/A vssd1 vssd1 vccd1 vccd1 _13581_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_197_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10792_ _15723_/Q _15789_/Q vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__and2b_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _11581_/B _15728_/Q vssd1 vssd1 vccd1 vccd1 _12531_/X sky130_fd_sc_hd__and2b_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13251__B _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15250_ _15347_/CLK _15250_/D _14299_/Y vssd1 vssd1 vccd1 vccd1 _15250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ _12462_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14201_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11987__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _15079_/Q _15244_/Q vssd1 vssd1 vccd1 vccd1 _11414_/C sky130_fd_sc_hd__and2_1
X_15181_ _15775_/CLK _15181_/D _14226_/Y vssd1 vssd1 vccd1 vccd1 _15181_/Q sky130_fd_sc_hd__dfrtp_1
X_12393_ _14943_/Q vssd1 vssd1 vccd1 vccd1 _12395_/A sky130_fd_sc_hd__inv_2
XANTENNA__14363__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14132_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1118 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11344_ _11344_/A _11344_/B vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__xor2_1
XFILLER_180_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08361__A _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14063_/Y sky130_fd_sc_hd__inv_2
X_11275_ _11275_/A _11275_/B _11275_/C vssd1 vssd1 vccd1 vccd1 _11277_/A sky130_fd_sc_hd__and3_1
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ _12945_/A _12944_/B _12942_/Y vssd1 vssd1 vccd1 vccd1 _13069_/B sky130_fd_sc_hd__a21o_1
X_10226_ _10225_/A _10225_/C _11402_/A vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _15147_/Q _15312_/Q vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14965_ _15727_/CLK _14965_/D _13997_/Y vssd1 vssd1 vccd1 vccd1 _14965_/Q sky130_fd_sc_hd__dfrtp_1
X_10088_ _10087_/A _10087_/B _10430_/A vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_output416_A _15589_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__A _15755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ input2/X vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__buf_6
XFILLER_48_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14896_ _15694_/CLK _14896_/D _13925_/Y vssd1 vssd1 vccd1 vccd1 _14896_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13847_ _13847_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13848_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14538__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater566_A _10933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13778_ _14983_/Q _13774_/A _13774_/B _13858_/B _14982_/Q vssd1 vssd1 vccd1 vccd1
+ _13778_/X sky130_fd_sc_hd__o311a_1
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15517_ _15553_/CLK _15517_/D _14582_/Y vssd1 vssd1 vccd1 vccd1 _15517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12729_ _12728_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__and2b_1
XFILLER_176_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater733_A _15675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _15569_/CLK _15448_/D _14509_/Y vssd1 vssd1 vccd1 vccd1 _15448_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11897__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater900_A input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15379_ _15750_/CLK _15379_/D _14435_/Y vssd1 vssd1 vccd1 vccd1 _15379_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_157_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14273__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09940_ _09939_/A _09939_/B _09993_/A vssd1 vssd1 vccd1 vccd1 _09946_/B sky130_fd_sc_hd__a21o_1
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09871_ _15185_/Q _09869_/Y _09875_/B vssd1 vssd1 vccd1 vccd1 _14955_/D sky130_fd_sc_hd__o21a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _15329_/Q _15345_/Q vssd1 vssd1 vccd1 vccd1 _08824_/A sky130_fd_sc_hd__or2b_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ _15414_/Q _07704_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__mux2_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _13145_/A _12970_/A vssd1 vssd1 vccd1 vccd1 _12667_/C sky130_fd_sc_hd__xor2_2
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07635_ _07635_/A vssd1 vssd1 vccd1 vccd1 _15448_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14448__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13352__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07566_ _07566_/A vssd1 vssd1 vccd1 vccd1 _15482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09305_ _15403_/Q _15387_/Q _09301_/B vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__o21a_1
XFILLER_210_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07497_ _07497_/A vssd1 vssd1 vccd1 vccd1 _15516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _15240_/D sky130_fd_sc_hd__xor2_2
XFILLER_166_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _15567_/Q _15547_/Q vssd1 vssd1 vccd1 vccd1 _09645_/A sky130_fd_sc_hd__xnor2_2
XFILLER_194_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_920 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14183__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ _08118_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__xnor2_1
XFILLER_79_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _15499_/Q _15483_/Q _09094_/B vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12415__B _12415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08049_ _11584_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11060_ _11052_/Y _11056_/B _11054_/B vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10011_ _15202_/Q _15103_/Q vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__or2b_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input147_A x_r_1[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/A vssd1 vssd1 vccd1 vccd1 _14750_/Y sky130_fd_sc_hd__inv_2
X_11962_ _12122_/A _11663_/C _11961_/Y vssd1 vssd1 vccd1 vccd1 _11963_/C sky130_fd_sc_hd__a21oi_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08678__A1 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13694_/A _13694_/B _13700_/X vssd1 vssd1 vccd1 vccd1 _13704_/A sky130_fd_sc_hd__o21ai_2
XFILLER_204_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ _14963_/Q _14897_/Q vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__or2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14681_/A vssd1 vssd1 vccd1 vccd1 _14681_/Y sky130_fd_sc_hd__inv_2
X_11893_ _11808_/A _11808_/B _11892_/X vssd1 vssd1 vccd1 vccd1 _11894_/B sky130_fd_sc_hd__a21oi_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14358__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ _09061_/A _13631_/B _09061_/B vssd1 vssd1 vccd1 vccd1 _15102_/D sky130_fd_sc_hd__a21boi_1
XFILLER_189_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844_ _10843_/A _10843_/C _10843_/B vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13563_ _15766_/Q _13563_/B vssd1 vssd1 vccd1 vccd1 _13564_/A sky130_fd_sc_hd__and2_1
XFILLER_158_725 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ _15720_/Q _15786_/Q vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12631__C1 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15302_ _15592_/CLK _15302_/D _14354_/Y vssd1 vssd1 vccd1 vccd1 _15302_/Q sky130_fd_sc_hd__dfrtp_1
X_12514_ _14953_/Q _12620_/B vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__xor2_1
XFILLER_13_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13494_/A _13782_/B vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__xor2_1
XFILLER_40_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15233_ _15700_/CLK _15233_/D _14282_/Y vssd1 vssd1 vccd1 vccd1 _15233_/Q sky130_fd_sc_hd__dfrtp_1
X_12445_ _12443_/Y _12445_/B vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__nand2b_1
XFILLER_139_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14093__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__A1 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15164_ _15729_/CLK _15164_/D _14208_/Y vssd1 vssd1 vccd1 vccd1 _15164_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08091__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _14941_/Q _12583_/B vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__and2_1
Xoutput509 output509/A vssd1 vssd1 vccd1 vccd1 y_r_6[4] sky130_fd_sc_hd__buf_2
XFILLER_153_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output366_A output366/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14115_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ _11327_/A _11327_/B _11327_/C vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__and3_1
XFILLER_158_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15095_ _15754_/CLK _15095_/D _14135_/Y vssd1 vssd1 vccd1 vccd1 _15095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14821__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14046_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14046_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11258_ _15778_/Q _15712_/Q vssd1 vssd1 vccd1 vccd1 _11259_/C sky130_fd_sc_hd__or2b_1
X_10209_ _10207_/Y _10209_/B vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13437__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__C _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11189_ _11365_/A _11190_/B vssd1 vssd1 vccd1 vccd1 _11189_/X sky130_fd_sc_hd__xor2_4
XFILLER_209_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater683_A _14488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _15790_/CLK _14948_/D _13980_/Y vssd1 vssd1 vccd1 vccd1 _14948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12995__B _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater850_A repeater851/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14879_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14268__A _14269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater948_A input150/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15802__D _15802_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07420_ _15553_/Q _07420_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _09021_/A _13614_/A vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__or2_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13111__S _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14731__A _14740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09923_ _09990_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__nand2_2
XFILLER_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _15753_/D sky130_fd_sc_hd__nor2_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _13895_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _15078_/D sky130_fd_sc_hd__xor2_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _15434_/Q _15418_/Q _09784_/X vssd1 vssd1 vccd1 vccd1 _09786_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ _08731_/X _08732_/Y _08734_/Y _08735_/X vssd1 vssd1 vccd1 vccd1 _08736_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_72_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_867 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08667_ _08728_/B _08433_/B _08666_/X vssd1 vssd1 vccd1 vccd1 _12658_/B sky130_fd_sc_hd__a21bo_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14178__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _15456_/Q input5/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07619_/A sky130_fd_sc_hd__mux2_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08598_/A _08598_/B vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__xor2_1
XFILLER_183_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07549_ _15490_/Q _07549_/A1 _07579_/S vssd1 vssd1 vccd1 vccd1 _07550_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_87_clk_A clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10558_/X _10565_/B vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__and2b_1
XFILLER_210_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08904__A _15456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_130_clk_A _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _15493_/Q _09219_/B _09219_/C vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__nand3_1
XFILLER_194_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10491_ _10963_/A _15284_/Q _10590_/B vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12230_ _12231_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_10_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12161_ _12161_/A _12117_/A vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__or2b_1
XFILLER_135_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14641__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11112_ _10877_/Y _11111_/B _10879_/B vssd1 vssd1 vccd1 vccd1 _11113_/B sky130_fd_sc_hd__o21ai_1
XFILLER_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12092_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _14927_/Q _14993_/Q vssd1 vssd1 vccd1 vccd1 _11044_/B sky130_fd_sc_hd__nand2_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07571__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__buf_12
XFILLER_18_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15782_ _15782_/CLK _15782_/D _14861_/Y vssd1 vssd1 vccd1 vccd1 _15782_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _13352_/A _13366_/A vssd1 vssd1 vccd1 vccd1 _12995_/C sky130_fd_sc_hd__xor2_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14733_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14733_/Y sky130_fd_sc_hd__inv_2
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ _11945_/A _11945_/B _12547_/A vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__or3_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14088__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14681_/A vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__inv_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11901_/B sky130_fd_sc_hd__nand2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13615_ _13614_/A _13614_/C _13614_/B vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__o21a_1
X_10827_ _15141_/Q _10826_/Y _10825_/B vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14595_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14595_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14816__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ _13546_/A _13546_/B vssd1 vssd1 vccd1 vccd1 _13547_/B sky130_fd_sc_hd__nand2_1
X_10758_ _11275_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10758_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_125_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output483_A _15621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13477_ _15771_/Q _13477_/B vssd1 vssd1 vccd1 vccd1 _13478_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _10689_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _11008_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__A _15757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15216_ _15347_/CLK _15216_/D _14264_/Y vssd1 vssd1 vccd1 vccd1 _15216_/Q sky130_fd_sc_hd__dfrtp_1
X_12428_ _12428_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _12455_/B sky130_fd_sc_hd__or2_1
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput306 output306/A vssd1 vssd1 vccd1 vccd1 y_i_2[5] sky130_fd_sc_hd__buf_2
Xoutput317 output317/A vssd1 vssd1 vccd1 vccd1 y_i_3[15] sky130_fd_sc_hd__buf_2
X_15147_ _15394_/CLK _15147_/D _14190_/Y vssd1 vssd1 vccd1 vccd1 _15147_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput328 output328/A vssd1 vssd1 vccd1 vccd1 y_i_4[0] sky130_fd_sc_hd__buf_2
X_12359_ _12357_/A _12575_/B _12358_/X vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__o21ai_1
Xoutput339 _11313_/Y vssd1 vssd1 vccd1 vccd1 y_i_4[4] sky130_fd_sc_hd__buf_2
XANTENNA__14551__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07864__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ _15758_/CLK _15078_/D _14117_/Y vssd1 vssd1 vccd1 vccd1 _15078_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater898_A input223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14029_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14029_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _09786_/A _09567_/B _09569_/X vssd1 vssd1 vccd1 vccd1 _09571_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ _12780_/A vssd1 vssd1 vccd1 vccd1 _08603_/B sky130_fd_sc_hd__inv_2
XFILLER_64_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12989__A3 _12976_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ _13012_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08455_/A sky130_fd_sc_hd__and2_1
XFILLER_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ _07403_/A vssd1 vssd1 vccd1 vccd1 _15566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08383_ _08411_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08412_/A sky130_fd_sc_hd__xor2_1
XFILLER_91_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14726__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12246__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _15371_/Q _15355_/Q vssd1 vssd1 vccd1 vccd1 _09005_/B sky130_fd_sc_hd__nand2_1
XFILLER_164_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__A2 _15420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _14960_/D sky130_fd_sc_hd__nor2_1
XFILLER_63_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09837_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _15749_/D sky130_fd_sc_hd__xor2_2
XFILLER_58_244 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07553__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13805__A _14986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ _15068_/Q _15101_/Q vssd1 vssd1 vccd1 vccd1 _09768_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08631_/X _08633_/A _08715_/Y _08717_/X _08718_/X vssd1 vssd1 vccd1 vccd1
+ _08719_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13524__B _13524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _15057_/Q _15090_/Q vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__nor2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11730_/A _11706_/A vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__or2b_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11661_ _11797_/A _11591_/B _11595_/B _11594_/X vssd1 vssd1 vccd1 vccd1 _11676_/A
+ sky130_fd_sc_hd__o31ai_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14636__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ _13769_/A _13400_/B vssd1 vssd1 vccd1 vccd1 _13747_/B sky130_fd_sc_hd__nand2_2
XFILLER_70_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10612_ _10612_/A _10612_/B _10612_/C vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__nor3_1
X_14380_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14399_/A sky130_fd_sc_hd__buf_12
XFILLER_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11592_ _11523_/A _11523_/B _11797_/A _08009_/C vssd1 vssd1 vccd1 vccd1 _11595_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13230_/A _13230_/B _13330_/Y vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__a21oi_1
XFILLER_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10543_ _10543_/A _10606_/A _10543_/C vssd1 vssd1 vccd1 vccd1 _10545_/A sky130_fd_sc_hd__or3_1
XFILLER_182_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input75_A x_i_4[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ _13263_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _13264_/A sky130_fd_sc_hd__nor2_1
X_10474_ _10473_/A _10473_/C _10473_/B vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ _15509_/CLK _15001_/D _14035_/Y vssd1 vssd1 vccd1 vccd1 _15001_/Q sky130_fd_sc_hd__dfrtp_2
X_12213_ _12213_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _12214_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14371__A _14376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ _13083_/A _13083_/B _13192_/X vssd1 vssd1 vccd1 vccd1 _13195_/B sky130_fd_sc_hd__a21oi_1
XFILLER_68_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09143__B_N _15562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _12144_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__or2_1
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _12075_/A _12075_/B _12075_/C vssd1 vssd1 vccd1 vccd1 _12186_/A sky130_fd_sc_hd__or3_1
XFILLER_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater809 _15578_/Q vssd1 vssd1 vccd1 vccd1 output421/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11026_ _11026_/A _11303_/B vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12977_ _13690_/A _13690_/B vssd1 vssd1 vccd1 vccd1 _13681_/B sky130_fd_sc_hd__nor2_2
X_15765_ _15774_/CLK _15765_/D _14844_/Y vssd1 vssd1 vccd1 vccd1 _15765_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11928_ _11928_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _11929_/B sky130_fd_sc_hd__nor2_1
X_14716_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14716_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13153__C _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15696_ _15768_/CLK _15696_/D _14771_/Y vssd1 vssd1 vccd1 vccd1 _15696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14647_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14647_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11859_ _11859_/A _11859_/B _11859_/C vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater646_A _11353_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14546__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_892 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14578_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14578_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13529_ _15759_/Q _13529_/B vssd1 vssd1 vccd1 vccd1 _13532_/C sky130_fd_sc_hd__nand2_1
XFILLER_201_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater813_A _15560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12066__A _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14281__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07594__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07783__A1 _07783_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ _10102_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__and2_1
XFILLER_29_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07883_ _07883_/A vssd1 vssd1 vccd1 vccd1 _15326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11844__S _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_1029 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09622_ _09621_/Y _15427_/Q _09617_/B vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__a21oi_1
XFILLER_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13608__A1 _15372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09553_ _15433_/Q _15417_/Q vssd1 vssd1 vccd1 vccd1 _09554_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13344__B _13746_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__xnor2_1
X_09484_ _09484_/A _09484_/B _09532_/A vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__nor3_1
XANTENNA__08157__C _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__xor2_1
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14456__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07769__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ _08366_/A _08384_/C vssd1 vssd1 vccd1 vccd1 _08376_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08454__A _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08297_ _11447_/C _08177_/Y _08296_/Y vssd1 vssd1 vccd1 vccd1 _08297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_558 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14191__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10190_ _10197_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13519__B _13519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10293__B_N _15153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07526__A1 _07526_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12900_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _12900_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_19_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _13880_/A _13880_/B vssd1 vssd1 vccd1 vccd1 _15056_/D sky130_fd_sc_hd__xnor2_1
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input227_A x_r_6[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ _12832_/A _12832_/B _12832_/C vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__a21o_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15571_/CLK _15550_/D _14616_/Y vssd1 vssd1 vccd1 vccd1 _15550_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _08583_/A _08583_/B _08700_/B _12691_/A _12692_/X vssd1 vssd1 vccd1 vccd1
+ _13057_/B sky130_fd_sc_hd__a311o_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14501_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14515_/A sky130_fd_sc_hd__buf_8
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11866_/A _11865_/C _11866_/B _11646_/A _11712_/X vssd1 vssd1 vccd1 vccd1
+ _11714_/B sky130_fd_sc_hd__a41o_1
XFILLER_159_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15525_/CLK _15481_/D _14544_/Y vssd1 vssd1 vccd1 vccd1 _15481_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12693_ _08583_/A _08583_/B _08700_/B _12692_/X vssd1 vssd1 vccd1 vccd1 _12694_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14366__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14432_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14432_/Y sky130_fd_sc_hd__inv_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11644_/A vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__inv_2
XFILLER_52_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14363_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14363_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11575_ _12369_/B _12369_/C _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11576_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 x_i_0[7] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput27 x_i_1[2] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13314_ _13273_/A _13273_/B _13272_/B vssd1 vssd1 vccd1 vccd1 _13315_/B sky130_fd_sc_hd__a21oi_2
Xinput38 x_i_2[12] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 x_i_2[8] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
X_10526_ _15258_/Q _15291_/Q vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14294_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output279_A output279/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13245_ _13244_/A _13244_/B _13244_/C vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_848 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10457_ _15125_/Q _10456_/Y _10455_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12889__A2 _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _13176_/A vssd1 vssd1 vccd1 vccd1 _13177_/B sky130_fd_sc_hd__inv_2
XFILLER_42_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10388_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _14941_/D sky130_fd_sc_hd__xor2_2
XANTENNA__07765__A1 input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output446_A _11369_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12127_ _12127_/A _12127_/B vssd1 vssd1 vccd1 vccd1 _12128_/B sky130_fd_sc_hd__nor2_2
XFILLER_123_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater606 _11363_/Y vssd1 vssd1 vccd1 vccd1 output443/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12058_ _12127_/A _12126_/C vssd1 vssd1 vccd1 vccd1 _12059_/B sky130_fd_sc_hd__or2b_1
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater617 _11169_/Y vssd1 vssd1 vccd1 vccd1 output509/A sky130_fd_sc_hd__clkbuf_2
Xrepeater628 _11161_/X vssd1 vssd1 vccd1 vccd1 output508/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater596_A _11183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater639 _10728_/Y vssd1 vssd1 vccd1 vccd1 output405/A sky130_fd_sc_hd__buf_4
X_11009_ _11008_/A _11008_/B _10689_/B vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08539__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15817_ _15817_/A vssd1 vssd1 vccd1 vccd1 _15817_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_repeater763_A _15639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15749_/CLK _15748_/D _14826_/Y vssd1 vssd1 vccd1 vccd1 _15748_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater930_A input173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15679_ _15679_/CLK _15679_/D _14753_/Y vssd1 vssd1 vccd1 vccd1 _15679_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14276__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08220_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08220_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__S _07589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_929 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_801 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08151_ _12254_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08082_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ _08986_/B _08984_/B vssd1 vssd1 vccd1 vccd1 _15103_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _11392_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__and2_1
XFILLER_25_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_704 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07508__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__A _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _15334_/Q _07866_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09605_ _09604_/A _09604_/B _09803_/A vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13074__B _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ _15368_/Q input236/X _07803_/S vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08168__B _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09536_ _09489_/A _09535_/B _09489_/B vssd1 vssd1 vccd1 vccd1 _15267_/D sky130_fd_sc_hd__a21boi_1
XFILLER_58_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _09466_/A _09466_/B _09522_/A vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14186__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08418_ _08418_/A _08645_/C vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08184__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _09398_/A _09398_/B _09398_/C vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__and3_1
XFILLER_200_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08349_ _12574_/B _12574_/C vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11360_ _11163_/Y _11359_/B _11165_/B vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__o21ai_2
XFILLER_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08912__A _08968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10311_ _10445_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _15779_/D sky130_fd_sc_hd__xnor2_4
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11291_ _15720_/Q _11290_/Y _11289_/B vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input177_A x_r_2[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ _13145_/A _13046_/A _13030_/C vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__and3_1
X_10242_ _15078_/Q _15243_/Q vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__or2_1
XFILLER_69_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11543__A2 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12740__A1 _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _15149_/Q _15314_/Q vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__and2b_1
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11992__B _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A x_i_2[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14981_ _15773_/CLK _14981_/D _14014_/Y vssd1 vssd1 vccd1 vccd1 _14981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13932_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13863_ _13863_/A _13863_/B _13863_/C vssd1 vssd1 vccd1 vccd1 _13865_/A sky130_fd_sc_hd__nor3_1
XFILLER_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ _12945_/A _12708_/X _12930_/A _12813_/X vssd1 vssd1 vccd1 vccd1 _12883_/B
+ sky130_fd_sc_hd__a31o_1
X_15602_ _15768_/CLK _15602_/D _14672_/Y vssd1 vssd1 vccd1 vccd1 _15602_/Q sky130_fd_sc_hd__dfrtp_2
X_13794_ _13794_/A _13801_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__xnor2_2
XFILLER_203_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12745_ _13145_/A _13319_/A vssd1 vssd1 vccd1 vccd1 _12784_/C sky130_fd_sc_hd__xor2_2
X_15533_ _15539_/CLK _15533_/D _14598_/Y vssd1 vssd1 vccd1 vccd1 _15533_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15630__D _15630_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14096__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_554 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07683__A0 _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ _15464_/CLK _15464_/D _14526_/Y vssd1 vssd1 vccd1 vccd1 _15464_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A _13037_/B vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__xnor2_1
XFILLER_175_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output396_A output396/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14415_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14415_/Y sky130_fd_sc_hd__inv_2
X_11627_ _11627_/A _11627_/B vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__xnor2_1
XFILLER_198_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15395_ _15575_/CLK _15395_/D _14453_/Y vssd1 vssd1 vccd1 vccd1 _15395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14346_/Y sky130_fd_sc_hd__inv_2
X_11558_ _11558_/A _11558_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__xor2_1
XFILLER_155_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10509_ _15287_/Q _15254_/Q vssd1 vssd1 vccd1 vccd1 _10510_/C sky130_fd_sc_hd__or2b_1
XANTENNA__09637__B _15544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14277_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14277_/Y sky130_fd_sc_hd__inv_2
X_11489_ _11489_/A _11542_/A vssd1 vssd1 vccd1 vccd1 _11491_/B sky130_fd_sc_hd__xnor2_1
XFILLER_171_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater609_A _11175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13228_ _13227_/B _12953_/C _13324_/A vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__o21ba_1
XFILLER_170_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__A1 _07738_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _13159_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13160_/B sky130_fd_sc_hd__and2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07872__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater880_A input247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater978_A repeater979/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _15406_/Q _07720_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07651_ _15440_/Q _07651_/A1 _07687_/S vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _07582_/A vssd1 vssd1 vccd1 vccd1 _15474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _09321_/A _09382_/A _09321_/C vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__nor3_1
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_913 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09252_ _09250_/X _09254_/C vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _12144_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _15569_/Q _15549_/Q _09182_/X vssd1 vssd1 vccd1 vccd1 _09188_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14734__A _14741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08134_ _15004_/Q vssd1 vssd1 vccd1 vccd1 _08223_/B sky130_fd_sc_hd__buf_6
XFILLER_175_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ _08066_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08118_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12254__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_976 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput206 x_r_4[5] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__clkbuf_2
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__A _15435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 x_r_5[15] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__clkbuf_1
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _08967_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _15197_/D sky130_fd_sc_hd__xor2_1
Xinput228 x_r_6[10] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput239 x_r_6[6] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__clkbuf_2
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ _09495_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__and2_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08898_ _15471_/Q _15455_/Q vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__or2b_1
XFILLER_5_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater970 repeater971/X vssd1 vssd1 vccd1 vccd1 _07386_/A1 sky130_fd_sc_hd__buf_4
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater981 input113/X vssd1 vssd1 vccd1 vccd1 repeater981/X sky130_fd_sc_hd__buf_2
X_07849_ _07849_/A vssd1 vssd1 vccd1 vccd1 _15343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10860_ _15775_/Q _11105_/B vssd1 vssd1 vccd1 vccd1 _10860_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _09518_/A _09518_/C _09518_/B vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__o21a_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10791_ _15722_/Q _15788_/Q vssd1 vssd1 vccd1 vccd1 _10795_/B sky130_fd_sc_hd__nand2_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _15728_/Q _11581_/B vssd1 vssd1 vccd1 vccd1 _12530_/X sky130_fd_sc_hd__or2b_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13251__C _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12461_ _12461_/A _12460_/Y vssd1 vssd1 vccd1 vccd1 _12462_/A sky130_fd_sc_hd__or2b_1
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14644__A _14661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14200_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__inv_2
X_11412_ _11412_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _15736_/D sky130_fd_sc_hd__nor2_2
X_15180_ _15180_/CLK _15180_/D _14225_/Y vssd1 vssd1 vccd1 vccd1 _15180_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11987__B _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12391_/A _12391_/C _12391_/B vssd1 vssd1 vccd1 vccd1 _12401_/C sky130_fd_sc_hd__a21o_1
XFILLER_165_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14131_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11343_ _14932_/Q _11342_/Y _11341_/B vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__a21o_1
XFILLER_193_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_818 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14062_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11274_ _15782_/Q _15716_/Q vssd1 vssd1 vccd1 vccd1 _11275_/C sky130_fd_sc_hd__or2b_1
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _13097_/B _13013_/B vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10225_ _10225_/A _11402_/A _10225_/C vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__and3_1
XFILLER_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _15146_/Q _15311_/Q vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__nand2_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14964_ _15777_/CLK _14964_/D _13996_/Y vssd1 vssd1 vccd1 vccd1 _14964_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10087_ _10087_/A _10087_/B _10430_/A vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__and3_1
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13521__B1_N _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13915_ _08841_/A _13914_/B _08841_/B vssd1 vssd1 vccd1 vccd1 _15069_/D sky130_fd_sc_hd__a21boi_1
XANTENNA_output311_A output311/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ _15383_/CLK _14895_/D _13924_/Y vssd1 vssd1 vccd1 vccd1 _14895_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10131__B _15307_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_684 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14819__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output409_A output409/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13846_ _14980_/Q _13846_/B vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__nand2_1
XFILLER_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13777_ _13860_/A _13777_/B vssd1 vssd1 vccd1 vccd1 _15705_/D sky130_fd_sc_hd__xnor2_1
XFILLER_90_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _15175_/Q _15274_/Q vssd1 vssd1 vccd1 vccd1 _10990_/C sky130_fd_sc_hd__or2b_1
XFILLER_15_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15516_ _15558_/CLK _15516_/D _14580_/Y vssd1 vssd1 vccd1 vccd1 _15516_/Q sky130_fd_sc_hd__dfrtp_2
X_12728_ _12729_/B _12728_/B vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__and2b_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12659_ _08671_/A _08671_/B _12658_/X vssd1 vssd1 vccd1 vccd1 _12768_/B sky130_fd_sc_hd__a21o_2
X_15447_ _15558_/CLK _15447_/D _14508_/Y vssd1 vssd1 vccd1 vccd1 _15447_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_repeater726_A _15690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14554__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07408__A0 _15563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15378_ _15724_/CLK _15378_/D _14434_/Y vssd1 vssd1 vccd1 vccd1 _15378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14329_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14329_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09870_ _10380_/A _15218_/Q _09971_/B vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__a21o_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A vssd1 vssd1 vccd1 vccd1 _15080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _13636_/A _13636_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10322__A _15126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ _07703_/A vssd1 vssd1 vccd1 vccd1 _15415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08683_ _13046_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__nand2_1
XFILLER_94_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14729__A _14739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A_N _15307_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _15448_/Q input12/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07635_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13352__B _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07565_ _15482_/Q _07565_/A1 _07579_/S vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09304_ _09302_/Y _09304_/B vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__nand2b_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07496_ _15516_/Q _07496_/A1 _07536_/S vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09235_ _09233_/A _09233_/B _09234_/X vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14464__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07777__S _07791_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09166_ _09642_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _15289_/D sky130_fd_sc_hd__xor2_1
XFILLER_119_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ _08290_/B vssd1 vssd1 vccd1 vccd1 _08118_/A sky130_fd_sc_hd__clkinv_4
XFILLER_163_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _09095_/Y _09097_/B vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__08181__B _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__A2 _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _08068_/A sky130_fd_sc_hd__xnor2_2
XFILLER_163_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_22 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12712__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10010_ _15103_/Q _15202_/Q vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__or2b_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08436__B1_N _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _09997_/A _09997_/B _09998_/X vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _12178_/A _12122_/A vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__nor2_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14639__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _10912_/A _10912_/B vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__nor2_1
X_13700_ _13700_/A _13700_/B vssd1 vssd1 vccd1 vccd1 _13700_/X sky130_fd_sc_hd__or2_1
XFILLER_56_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14680_/A vssd1 vssd1 vccd1 vccd1 _14680_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11892_ _11892_/A _11892_/B vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__and2_1
XFILLER_204_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ _13631_/A _13631_/B vssd1 vssd1 vccd1 vccd1 _15101_/D sky130_fd_sc_hd__xnor2_1
X_10843_ _10843_/A _10843_/B _10843_/C vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__and3_1
XANTENNA__09627__A1 _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07638__A0 _15446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13562_ _13564_/B _13562_/B vssd1 vssd1 vccd1 vccd1 _15602_/D sky130_fd_sc_hd__nor2_1
XFILLER_73_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10774_ _10774_/A _11287_/B vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__nand2_1
XFILLER_198_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12513_ _12520_/A _12520_/B vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__xnor2_2
XFILLER_158_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15301_ _15592_/CLK _15301_/D _14353_/Y vssd1 vssd1 vccd1 vccd1 _15301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _13790_/A _13790_/B vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14374__A _14379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07687__S _07687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ _12444_/A _12463_/B _12463_/C vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__nand3_1
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15232_ _15506_/CLK _15232_/D _14281_/Y vssd1 vssd1 vccd1 vccd1 _15232_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08372__A _08396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11737__A2 _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15163_ _15699_/CLK _15163_/D _14207_/Y vssd1 vssd1 vccd1 vccd1 _15163_/Q sky130_fd_sc_hd__dfrtp_1
X_12375_ _12375_/A _12582_/A vssd1 vssd1 vccd1 vccd1 _15646_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14114_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _14994_/Q _14928_/Q vssd1 vssd1 vccd1 vccd1 _11327_/C sky130_fd_sc_hd__or2b_1
XFILLER_153_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15094_ _15110_/CLK _15094_/D _14134_/Y vssd1 vssd1 vccd1 vccd1 _15094_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output261_A output261/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output359_A _15683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14045_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11259_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10208_ _15073_/Q _15238_/Q vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__nand2_1
X_11188_ _15748_/Q _11187_/Y _11183_/B vssd1 vssd1 vccd1 vccd1 _11190_/B sky130_fd_sc_hd__a21o_1
XANTENNA_output526_A output526/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__B1 _11369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11238__A _15034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _10832_/A _10139_/B vssd1 vssd1 vccd1 vccd1 _15800_/D sky130_fd_sc_hd__xor2_1
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14947_ _15790_/CLK _14947_/D _13979_/Y vssd1 vssd1 vccd1 vccd1 _14947_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater676_A _14559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14549__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13453__A _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14878_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14878_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13829_ _13829_/A _13829_/B vssd1 vssd1 vccd1 vccd1 _15667_/D sky130_fd_sc_hd__xnor2_4
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14284__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ _15374_/Q _15358_/Q vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__and2_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10317__A _15125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _15194_/Q _15227_/Q vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09853_ _09852_/A _09852_/C _09852_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__a21oi_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _13893_/A _08798_/B _08803_/X vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__a21o_1
X_09784_ _15434_/Q _15418_/Q _09783_/B vssd1 vssd1 vccd1 vccd1 _09784_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08735_ _12881_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _08735_/X sky130_fd_sc_hd__or2_1
XFILLER_67_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14459__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__A0 _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11664__A1 _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08666_ _08666_/A _08432_/A vssd1 vssd1 vccd1 vccd1 _08666_/X sky130_fd_sc_hd__or2b_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07617_ _07617_/A vssd1 vssd1 vccd1 vccd1 _15457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _08597_/A _08621_/A vssd1 vssd1 vccd1 vccd1 _08598_/B sky130_fd_sc_hd__nand2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07548_ _07548_/A vssd1 vssd1 vccd1 vccd1 _15491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14194__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _15524_/Q _07479_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12707__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _15493_/Q _09219_/B _09219_/C vssd1 vssd1 vccd1 vccd1 _09222_/C sky130_fd_sc_hd__a21o_1
XFILLER_210_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ _15284_/Q _10590_/B vssd1 vssd1 vccd1 vccd1 _10490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12426__B _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09149_ _15563_/Q _15543_/Q vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__and2_1
XFILLER_33_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _12160_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__or2b_1
XFILLER_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11111_ _11111_/A _11111_/B vssd1 vssd1 vccd1 vccd1 _11111_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_190_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _12149_/A _12148_/C vssd1 vssd1 vccd1 vccd1 _12092_/B sky130_fd_sc_hd__or2b_1
XANTENNA_input257_A x_r_7[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_967 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _14927_/Q _14993_/Q vssd1 vssd1 vccd1 vccd1 _11042_/Y sky130_fd_sc_hd__nor2_1
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14801_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input20_A x_i_1[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15782_/CLK _15781_/D _14860_/Y vssd1 vssd1 vccd1 vccd1 _15781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14369__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ _12993_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13273__A _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14732_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14732_/Y sky130_fd_sc_hd__inv_2
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11944_ _12548_/A _12549_/A vssd1 vssd1 vccd1 vccd1 _12547_/A sky130_fd_sc_hd__nand2_2
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08367__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _15732_/Q _11875_/B vssd1 vssd1 vccd1 vccd1 _11945_/A sky130_fd_sc_hd__and2_1
X_14663_ _14675_/A vssd1 vssd1 vccd1 vccd1 _14663_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10826_ _15306_/Q vssd1 vssd1 vccd1 vccd1 _10826_/Y sky130_fd_sc_hd__inv_2
X_13614_ _13614_/A _13614_/B _13614_/C vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__nor3_1
XFILLER_38_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14594_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A2 _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _10751_/A _10753_/B _10751_/B vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__a21boi_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13545_ _13545_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__or2_1
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_clk clkbuf_opt_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15693_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11521__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13476_ _15771_/Q _13477_/B vssd1 vssd1 vccd1 vccd1 _13478_/A sky130_fd_sc_hd__or2_1
X_10688_ _15180_/Q _15279_/Q vssd1 vssd1 vccd1 vccd1 _10689_/B sky130_fd_sc_hd__and2b_1
XFILLER_139_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output476_A output476/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12427_ _12439_/B _12427_/B vssd1 vssd1 vccd1 vccd1 _12428_/B sky130_fd_sc_hd__and2_1
XFILLER_12_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15215_ _15347_/CLK _15215_/D _14263_/Y vssd1 vssd1 vccd1 vccd1 _15215_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14832__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput307 output307/A vssd1 vssd1 vccd1 vccd1 y_i_2[6] sky130_fd_sc_hd__buf_2
X_12358_ _12358_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12358_/X sky130_fd_sc_hd__or2_1
X_15146_ _15394_/CLK _15146_/D _14189_/Y vssd1 vssd1 vccd1 vccd1 _15146_/Q sky130_fd_sc_hd__dfrtp_2
Xoutput318 output318/A vssd1 vssd1 vccd1 vccd1 y_i_3[16] sky130_fd_sc_hd__buf_2
XFILLER_58_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput329 _11338_/X vssd1 vssd1 vccd1 vccd1 y_i_4[10] sky130_fd_sc_hd__buf_2
XFILLER_141_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15077_ _15754_/CLK _15077_/D _14116_/Y vssd1 vssd1 vccd1 vccd1 _15077_/Q sky130_fd_sc_hd__dfrtp_1
X_12289_ _12289_/A _12289_/B vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12352__A _14939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14028_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14028_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater793_A _15598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07880__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater960_A input134/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08520_ _12871_/A _12780_/A _08520_/C vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__and3_1
XFILLER_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ _08451_/A _08451_/B vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07402_ _15566_/Q input126/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__mux2_1
X_08382_ _13366_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_195_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_124_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15501_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11431__A _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09003_ _15371_/Q _15355_/Q vssd1 vssd1 vccd1 vccd1 _09003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12262__A _12262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__B _15416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _09904_/A _09904_/C _09981_/A vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__a21oi_1
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09836_ _15059_/Q _09835_/Y _09834_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__a21o_1
XFILLER_98_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _09767_/A _09863_/A vssd1 vssd1 vccd1 vccd1 _15724_/D sky130_fd_sc_hd__xor2_2
XANTENNA__14189__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15723__D _15723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08718_ _08718_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _08718_/X sky130_fd_sc_hd__or2_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09822_/A _09698_/B vssd1 vssd1 vccd1 vccd1 _15712_/D sky130_fd_sc_hd__xnor2_1
XFILLER_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08187__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08649_/A _08649_/B vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__xnor2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11607_/A _11607_/B _11659_/X vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__a21o_1
XFILLER_25_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ _15261_/Q _15294_/Q vssd1 vssd1 vccd1 vccd1 _10612_/C sky130_fd_sc_hd__and2_1
XFILLER_211_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _11797_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_115_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15700_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13032__S _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _13330_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10542_ _15292_/Q _15259_/Q vssd1 vssd1 vccd1 vccd1 _10543_/C sky130_fd_sc_hd__and2b_1
XFILLER_183_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_576 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ _13350_/A _13261_/B vssd1 vssd1 vccd1 vccd1 _13263_/B sky130_fd_sc_hd__and2_1
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _10473_/A _10473_/B _10473_/C vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__and3_1
XFILLER_183_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14652__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _12213_/A _12482_/A vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__and2_1
XFILLER_170_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15000_ _15509_/CLK _15000_/D _14034_/Y vssd1 vssd1 vccd1 vccd1 _15000_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _13082_/B _13192_/B vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__and2b_1
XFILLER_136_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input68_A x_i_4[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12143_ _12144_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13314__A1 _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _12074_/A _12074_/B vssd1 vssd1 vccd1 vccd1 _12075_/C sky130_fd_sc_hd__xnor2_1
XFILLER_151_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11025_ _11023_/Y _11025_/B vssd1 vssd1 vccd1 vccd1 _11303_/B sky130_fd_sc_hd__and2b_1
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14099__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/CLK _15764_/D _14843_/Y vssd1 vssd1 vccd1 vccd1 _15764_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08097__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _12976_/A _12976_/B _12976_/C vssd1 vssd1 vccd1 vccd1 _13690_/B sky130_fd_sc_hd__and3_1
XFILLER_45_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14715_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14715_/Y sky130_fd_sc_hd__inv_2
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11927_ _11928_/A _11928_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__and2_1
XFILLER_166_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15695_ _15775_/CLK _15695_/D _14770_/Y vssd1 vssd1 vccd1 vccd1 _15695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14646_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _11859_/A _11859_/B _11859_/C vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__a21o_1
XFILLER_177_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10809_ _10809_/A _10809_/B _10809_/C vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_106_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15770_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_repeater541_A _11296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _11789_/A _12540_/A vssd1 vssd1 vccd1 vccd1 _15582_/D sky130_fd_sc_hd__xor2_1
X_14577_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14577_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater639_A _10728_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13528_ _13530_/A _13528_/B vssd1 vssd1 vccd1 vccd1 _15595_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__12066__B _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_846 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater806_A _15583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13461_/C sky130_fd_sc_hd__xnor2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14562__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_71_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15808__D _15808_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13178__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15129_ _15433_/CLK _15129_/D _14171_/Y vssd1 vssd1 vccd1 vccd1 _15129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07951_ _15119_/Q _15284_/Q vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__or2_1
XFILLER_101_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_86_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _15326_/Q input146/X _07892_/S vssd1 vssd1 vccd1 vccd1 _07883_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12810__A _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _15443_/Q vssd1 vssd1 vccd1 vccd1 _09621_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_896 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13608__A2 _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09552_ _15433_/Q _15417_/Q vssd1 vssd1 vccd1 vccd1 _09552_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ _08508_/B _08503_/B vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _15539_/Q _15523_/Q vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14737__A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08434_ _08728_/B _08434_/B vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08735__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ _12921_/A _12810_/A vssd1 vssd1 vccd1 vccd1 _08384_/C sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_leaf_24_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08454__B _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08296_ _11435_/A _11467_/A _08295_/X vssd1 vssd1 vccd1 vccd1 _08296_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_192_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07471__A1 _07471_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _15044_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__14472__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08470__A _14907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09819_ _15088_/Q vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input122_A x_i_7[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ _12883_/B _12830_/B vssd1 vssd1 vccd1 vccd1 _12832_/C sky130_fd_sc_hd__xor2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12283__A1 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12807_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__xor2_2
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14647__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14500_/Y sky130_fd_sc_hd__inv_2
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11570_/A _11643_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11712_/X sky130_fd_sc_hd__o21a_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15480_ _15569_/CLK _15480_/D _14543_/Y vssd1 vssd1 vccd1 vccd1 _15480_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12692_ _08699_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__and2b_1
XFILLER_188_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08645__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11643_ _11643_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11644_/A sky130_fd_sc_hd__or2b_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__inv_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _11648_/A _11648_/B _12369_/B _12369_/C vssd1 vssd1 vccd1 vccd1 _11576_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_161_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_863 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09110__B_N _15503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14362_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14362_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 x_i_0[8] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput28 x_i_1[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
Xinput39 x_i_2[13] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13313_ _13369_/B _13313_/B vssd1 vssd1 vccd1 vccd1 _13315_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10525_ _15258_/Q _15291_/Q vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__or2_1
XFILLER_183_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14293_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14293_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14382__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13244_ _13244_/A _13244_/B _13244_/C vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__and3_1
XFILLER_183_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10456_ _15158_/Q vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11213__B_N _15031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__A _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13175_/A _13175_/B vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__or2_1
XFILLER_123_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10387_ _15203_/Q _10386_/Y _10385_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__a21o_1
X_12126_ _12126_/A _12126_/B _12126_/C vssd1 vssd1 vccd1 vccd1 _12127_/B sky130_fd_sc_hd__and3_1
XFILLER_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output341_A output341/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output439_A output439/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12057_ _12056_/A _12056_/B _12056_/C vssd1 vssd1 vccd1 vccd1 _12126_/C sky130_fd_sc_hd__a21o_1
XFILLER_133_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater607 _11316_/X vssd1 vssd1 vccd1 vccd1 output340/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12630__A _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater618 _11113_/Y vssd1 vssd1 vccd1 vccd1 output374/A sky130_fd_sc_hd__clkbuf_2
Xrepeater629 _11031_/Y vssd1 vssd1 vccd1 vccd1 output270/A sky130_fd_sc_hd__clkbuf_2
X_11008_ _11008_/A _11008_/B vssd1 vssd1 vccd1 vccd1 _15016_/D sky130_fd_sc_hd__xor2_1
XFILLER_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_896 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15816_ _15816_/A vssd1 vssd1 vccd1 vccd1 _15816_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12274__A1 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15749_/CLK _15747_/D _14825_/Y vssd1 vssd1 vccd1 vccd1 _15747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12959_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_repeater756_A _15646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14557__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15678_ _15679_/CLK _15678_/D _14752_/Y vssd1 vssd1 vccd1 vccd1 _15678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_988 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14629_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14629_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater923_A input186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _08150_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08081_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08081_/X sky130_fd_sc_hd__or2_1
XANTENNA__07453__A1 _07453_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14292__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08290__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A1 _15468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ _15365_/Q _08983_/B _13591_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__and3_1
XFILLER_102_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _15053_/Q _15218_/Q vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__or2_1
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_716 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _07865_/A vssd1 vssd1 vccd1 vccd1 _15335_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09604_/A _09604_/B _09803_/A vssd1 vssd1 vccd1 vccd1 _09604_/X sky130_fd_sc_hd__and3_1
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07796_ _07796_/A vssd1 vssd1 vccd1 vccd1 _15369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _15266_/D sky130_fd_sc_hd__xnor2_1
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14467__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _09466_/A _09466_/B _09522_/A vssd1 vssd1 vccd1 vccd1 _09466_/X sky130_fd_sc_hd__and3_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08417_ _13012_/A _12921_/A vssd1 vssd1 vccd1 vccd1 _08645_/C sky130_fd_sc_hd__xor2_1
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _09397_/A _09397_/B vssd1 vssd1 vccd1 vccd1 _09398_/C sky130_fd_sc_hd__nand2_1
XFILLER_71_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__A_N _15426_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08184__B _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _08347_/B _08347_/C _08347_/A vssd1 vssd1 vccd1 vccd1 _12574_/C sky130_fd_sc_hd__a21oi_1
XFILLER_132_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08279_ _08279_/A _08279_/B vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__xnor2_2
XFILLER_164_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12715__A _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10304_/A _10306_/B _10304_/B vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__a21boi_4
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11290_ _15786_/Q vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10241_ _10241_/A _10241_/B vssd1 vssd1 vccd1 vccd1 _15766_/D sky130_fd_sc_hd__nor2_1
XFILLER_154_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10172_ _15148_/Q _15313_/Q vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11765__S _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput490 _15612_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[2] sky130_fd_sc_hd__buf_2
XFILLER_105_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14980_ _15773_/CLK _14980_/D _14013_/Y vssd1 vssd1 vccd1 vccd1 _14980_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13931_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13931_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _14983_/Q _13862_/B vssd1 vssd1 vccd1 vccd1 _13863_/C sky130_fd_sc_hd__and2_1
XFILLER_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15601_ _15773_/CLK _15601_/D _14671_/Y vssd1 vssd1 vccd1 vccd1 _15601_/Q sky130_fd_sc_hd__dfrtp_1
X_12813_ _12640_/A _12813_/B _12813_/C vssd1 vssd1 vccd1 vccd1 _12813_/X sky130_fd_sc_hd__and3b_1
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13793_ _13785_/A _13785_/B _13792_/X vssd1 vssd1 vccd1 vccd1 _13801_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14377__A _14379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13281__A _13737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15532_ _15532_/CLK _15532_/D _14597_/Y vssd1 vssd1 vccd1 vccd1 _15532_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _13046_/A _13220_/A vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07683__A1 input181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11513__B _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15493_/CLK _15463_/D _14525_/Y vssd1 vssd1 vccd1 vccd1 _15463_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12675_ _13046_/A _13220_/A vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__xor2_2
X_14414_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14414_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11626_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15394_ _15394_/CLK _15394_/D _14452_/Y vssd1 vssd1 vccd1 vccd1 _15394_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output389_A _15695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07435__A1 _07435_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14345_/Y sky130_fd_sc_hd__inv_2
X_11557_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__xor2_1
XFILLER_155_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10508_ _10506_/Y _10508_/B vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__and2b_1
X_11488_ _08176_/A _08174_/X _08175_/A vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__a21oi_1
X_14276_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14276_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _14890_/D sky130_fd_sc_hd__nor2_1
X_13227_ _13438_/A _13227_/B vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__and2_1
XFILLER_48_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14840__A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _13159_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12178_/A _12122_/A vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__nand2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13089_ _13089_/A _13089_/B vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater873_A repeater874/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ _07650_/A vssd1 vssd1 vccd1 vccd1 _15441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _15474_/Q input71/X _07591_/S vssd1 vssd1 vccd1 vccd1 _07582_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14287__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09320_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _09321_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ _09250_/B _09250_/C _09250_/A vssd1 vssd1 vccd1 vccd1 _09254_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08399__C_N _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08202_ _12088_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09182_ _15569_/Q _15549_/Q _09178_/B vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08133_ _11491_/A _08223_/C vssd1 vssd1 vccd1 vccd1 _08236_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07426__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08064_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_988 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14750__A _14750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput207 x_r_4[6] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13366__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput218 x_r_5[1] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__clkbuf_2
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09563__B _15419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput229 x_r_6[11] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__clkbuf_2
X_08966_ _15472_/Q _15456_/Q _08965_/B vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07917_ _15525_/Q _15509_/Q vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__or2_1
XFILLER_97_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08897_ _15455_/Q _15471_/Q vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__or2b_1
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15374_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater960 input134/X vssd1 vssd1 vccd1 vccd1 _07876_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_17_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater971 input119/X vssd1 vssd1 vccd1 vccd1 repeater971/X sky130_fd_sc_hd__buf_2
X_07848_ _15343_/Q _07848_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater982 input112/X vssd1 vssd1 vccd1 vccd1 _07528_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14197__A _14198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07779_ _15377_/Q _07779_/A1 _07791_/S vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15731__D _15731_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ _09518_/A _09518_/B _09518_/C vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__nor3_1
X_10790_ _10790_/A vssd1 vssd1 vccd1 vccd1 _10790_/X sky130_fd_sc_hd__clkbuf_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07665__A1 _07665_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09449_ _09449_/A _09518_/A vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__or2_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_738 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ _12460_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ _11411_/A _11411_/B _11411_/C vssd1 vssd1 vccd1 vccd1 _11414_/B sky130_fd_sc_hd__and3_1
XFILLER_184_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12391_ _12391_/A _12391_/B _12391_/C vssd1 vssd1 vccd1 vccd1 _12401_/B sky130_fd_sc_hd__nand3_1
XFILLER_193_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_676 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14130_ _14138_/A vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11342_ _14998_/Q vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11273_ _11273_/A _11273_/B vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__nand2_1
X_14061_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14660__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input50_A x_i_2[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _13012_/A _13012_/B vssd1 vssd1 vccd1 vccd1 _13013_/B sky130_fd_sc_hd__or2_1
X_10224_ _15239_/Q _15074_/Q vssd1 vssd1 vccd1 vccd1 _10225_/C sky130_fd_sc_hd__or2b_1
XFILLER_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_906 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10155_ _10155_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14963_ _15775_/CLK _14963_/D _13995_/Y vssd1 vssd1 vccd1 vccd1 _14963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__nor2_2
XFILLER_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13914_ _13914_/A _13914_/B vssd1 vssd1 vccd1 vccd1 _15068_/D sky130_fd_sc_hd__xnor2_1
X_14894_ _15383_/CLK _14894_/D _13923_/Y vssd1 vssd1 vccd1 vccd1 _14894_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13845_ _13845_/A vssd1 vssd1 vccd1 vccd1 _15670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output304_A output304/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11524__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13776_ _13767_/A _13767_/B _13858_/B _14982_/Q vssd1 vssd1 vccd1 vccd1 _13777_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__nand2_1
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12339__B _12339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15515_ _15749_/CLK _15515_/D _14579_/Y vssd1 vssd1 vccd1 vccd1 _15515_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12727_ _12654_/A _12654_/B _12726_/X vssd1 vssd1 vccd1 vccd1 _12728_/B sky130_fd_sc_hd__a21bo_1
XFILLER_204_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14835__A _14836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15446_ _15511_/CLK _15446_/D _14507_/Y vssd1 vssd1 vccd1 vccd1 _15446_/Q sky130_fd_sc_hd__dfrtp_4
X_12658_ _08668_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07408__A1 _07408_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11609_ _11658_/A _11658_/B vssd1 vssd1 vccd1 vccd1 _11611_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_repeater621_A _10883_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15377_ _15724_/CLK _15377_/D _14433_/Y vssd1 vssd1 vccd1 vccd1 _15377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ _12395_/Y _12588_/B _12396_/A vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__a21oi_1
XFILLER_117_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater719_A _15700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14328_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14328_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14570__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08818_/X _08825_/B vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08751_ _08751_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _13636_/B sky130_fd_sc_hd__or2b_1
XFILLER_57_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _15717_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07702_ _15415_/Q _07702_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08682_ _14918_/Q vssd1 vssd1 vccd1 vccd1 _13491_/S sky130_fd_sc_hd__buf_4
XFILLER_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _07633_/A vssd1 vssd1 vccd1 vccd1 _15449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07564_ _07564_/A vssd1 vssd1 vccd1 vccd1 _15483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_560 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ _15404_/Q _15388_/Q vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07647__A1 _07647_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07495_ _07495_/A vssd1 vssd1 vccd1 vccd1 _15517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14745__A _14751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_587 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _15498_/Q _15482_/Q vssd1 vssd1 vccd1 vccd1 _09234_/X sky130_fd_sc_hd__and2b_1
XFILLER_210_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09165_ _15565_/Q _15545_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08116_ _08120_/C _08112_/A _08112_/B _08325_/A _08325_/B vssd1 vssd1 vccd1 vccd1
+ _08323_/B sky130_fd_sc_hd__a32o_1
XFILLER_108_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ _15500_/Q _15484_/Q vssd1 vssd1 vccd1 vccd1 _09097_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _08047_/A _11434_/A vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_162_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14480__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07793__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_34 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12712__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11609__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _15197_/Q _15230_/Q vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__and2_1
XFILLER_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ _15466_/Q _15450_/Q _08948_/X vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk _15666_/CLK vssd1 vssd1 vccd1 vccd1 _15688_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _11960_/A _12055_/A _11977_/A vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__and3_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _10910_/A _10910_/C _11119_/A vssd1 vssd1 vccd1 vccd1 _10912_/B sky130_fd_sc_hd__a21oi_1
Xrepeater790 _15602_/Q vssd1 vssd1 vccd1 vccd1 output462/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07886__A1 _07886_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11891_ _11891_/A _11891_/B vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__nand2_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13630_ _15379_/Q _15363_/Q _13629_/X vssd1 vssd1 vccd1 vccd1 _13631_/B sky130_fd_sc_hd__a21o_1
XANTENNA_input202_A x_r_4[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _10842_/A vssd1 vssd1 vccd1 vccd1 _14914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07638__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__A1 _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13561_ _13561_/A _13561_/B _13561_/C vssd1 vssd1 vccd1 vccd1 _13562_/B sky130_fd_sc_hd__and3_1
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10773_ _10774_/A _11287_/B vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__xor2_1
XANTENNA__14655__A _14656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15300_ _15563_/CLK _15300_/D _14352_/Y vssd1 vssd1 vccd1 vccd1 _15300_/Q sky130_fd_sc_hd__dfrtp_1
X_12512_ _12502_/A _12502_/B _12511_/Y vssd1 vssd1 vccd1 vccd1 _12520_/B sky130_fd_sc_hd__o21a_1
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input98_A x_i_5[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08653__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ _13492_/A _13492_/B vssd1 vssd1 vccd1 vccd1 _13790_/B sky130_fd_sc_hd__xnor2_4
XFILLER_201_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15231_ _15506_/CLK _15231_/D _14279_/Y vssd1 vssd1 vccd1 vccd1 _15231_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _12463_/B _12463_/C _12444_/A vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08372__B _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08063__A1 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ _15699_/CLK _15162_/D _14206_/Y vssd1 vssd1 vccd1 vccd1 _15162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12374_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__xnor2_2
XFILLER_158_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14113_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14113_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07810__A1 input167/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11327_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14390__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15750_/CLK _15093_/D _14133_/Y vssd1 vssd1 vccd1 vccd1 _15093_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14044_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11256_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__xor2_2
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11519__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _15073_/Q _15238_/Q vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__nor2_1
X_11187_ _15026_/Q vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11370__A1 _15751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _10132_/A _10134_/B _10132_/B vssd1 vssd1 vccd1 vccd1 _10139_/B sky130_fd_sc_hd__a21boi_1
XANTENNA_output421_A output421/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15729_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output519_A output519/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14946_ _15784_/CLK _14946_/D _13977_/Y vssd1 vssd1 vccd1 vccd1 _14946_/Q sky130_fd_sc_hd__dfrtp_1
X_10069_ _15114_/Q _15213_/Q vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__and2b_1
XFILLER_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14877_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14877_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater571_A repeater572/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater669_A _14709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13828_ _13696_/B _13826_/B _13827_/X vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__a21o_1
XFILLER_189_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13743_/A _13842_/A _13848_/A _13758_/X vssd1 vssd1 vccd1 vccd1 _13767_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_188_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater836_A input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14565__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07878__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15429_ _15808_/CLK _15429_/D _14489_/Y vssd1 vssd1 vccd1 vccd1 _15429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07801__A1 _07801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09921_ _15194_/Q _15227_/Q vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__or2_1
XANTENNA__07907__A _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08502__S _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09852_/A _09852_/B _09852_/C vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__and3_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08803_ _15341_/Q _15325_/Q vssd1 vssd1 vccd1 vccd1 _08803_/X sky130_fd_sc_hd__and2b_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09783_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _15157_/D sky130_fd_sc_hd__xnor2_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08734_ _12921_/A _12871_/A vssd1 vssd1 vccd1 vccd1 _08734_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_6_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__A1 input195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11664__A2 _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _12627_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _08668_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__15281__D _15281_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _15457_/Q _07616_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08596_ _08596_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _08718_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07547_ _15491_/Q input40/X _07579_/S vssd1 vssd1 vccd1 vccd1 _07548_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14475__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07478_ _07478_/A vssd1 vssd1 vccd1 vccd1 _15525_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08473__A _14908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09217_ _15477_/Q vssd1 vssd1 vccd1 vccd1 _09219_/B sky130_fd_sc_hd__inv_2
XFILLER_33_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09148_ _15562_/Q _15542_/Q _09147_/B vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__a21oi_1
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _15496_/Q _15480_/Q vssd1 vssd1 vccd1 vccd1 _09080_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11110_ _10872_/A _11109_/B _10872_/B vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__a21boi_1
XFILLER_135_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12090_ _12089_/A _12089_/B _12089_/C vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__a21o_1
XFILLER_122_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08348__A2 _08347_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11317_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input152_A x_r_1[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14800_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15780_ _15782_/CLK _15780_/D _14859_/Y vssd1 vssd1 vccd1 vccd1 _15780_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _12992_/A _12992_/B vssd1 vssd1 vccd1 vccd1 _13008_/B sky130_fd_sc_hd__or2_1
XFILLER_58_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14731_/Y sky130_fd_sc_hd__inv_2
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A x_i_0[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _15733_/Q _11950_/B vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__or2_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__buf_6
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _11874_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _15583_/D sky130_fd_sc_hd__nor2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _09021_/A _13613_/B vssd1 vssd1 vccd1 vccd1 _13614_/C sky130_fd_sc_hd__and2b_1
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _14910_/D sky130_fd_sc_hd__nor2_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14593_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14385__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08284__A1 _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ _13544_/A vssd1 vssd1 vccd1 vccd1 _15598_/D sky130_fd_sc_hd__clkbuf_1
X_10756_ _10754_/Y _10756_/B vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__and2b_1
XFILLER_197_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11521__B _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13475_ _13475_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13477_/B sky130_fd_sc_hd__xnor2_1
XFILLER_173_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10687_ _15279_/Q _15180_/Q vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__and2b_1
XFILLER_173_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15214_ _15347_/CLK _15214_/D _14262_/Y vssd1 vssd1 vccd1 vccd1 _15214_/Q sky130_fd_sc_hd__dfrtp_1
X_12426_ _11952_/B _12426_/B vssd1 vssd1 vccd1 vccd1 _12430_/C sky130_fd_sc_hd__and2b_1
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output371_A _11107_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output469_A output469/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput308 _10905_/X vssd1 vssd1 vccd1 vccd1 y_i_2[7] sky130_fd_sc_hd__buf_2
X_15145_ _15394_/CLK _15145_/D _14188_/Y vssd1 vssd1 vccd1 vccd1 _15145_/Q sky130_fd_sc_hd__dfrtp_1
X_12357_ _12357_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _15644_/D sky130_fd_sc_hd__xor2_1
XFILLER_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput319 _15661_/Q vssd1 vssd1 vccd1 vccd1 y_i_3[1] sky130_fd_sc_hd__buf_2
XANTENNA__07795__A0 _15369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12633__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08830__B _15330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11308_/X sky130_fd_sc_hd__xor2_4
X_15076_ _15249_/CLK _15076_/D _14115_/Y vssd1 vssd1 vccd1 vccd1 _15076_/Q sky130_fd_sc_hd__dfrtp_1
X_12288_ _12260_/A _12260_/B _12257_/A vssd1 vssd1 vccd1 vccd1 _12289_/B sky130_fd_sc_hd__a21oi_1
XFILLER_153_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14027_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14027_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11239_ _15756_/Q _11238_/Y _11237_/B vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__07547__A0 _15491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09942__A _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater786_A _15606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_931 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13183__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ _15501_/CLK _14929_/D _13960_/Y vssd1 vssd1 vccd1 vccd1 _14929_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater953_A input143/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _08459_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08451_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_986 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07401_ _07401_/A vssd1 vssd1 vccd1 vccd1 _15567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08381_ _08381_/A _08422_/C vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__xnor2_1
XFILLER_211_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14295__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08293__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10328__A _15127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09002_ _13602_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _15107_/D sky130_fd_sc_hd__xor2_1
XFILLER_118_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15276__D _15276_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _09904_/A _09981_/A _09904_/C vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__and3_1
XFILLER_99_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07538__A0 _15495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input5_A x_i_0[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _15092_/Q vssd1 vssd1 vccd1 vccd1 _09835_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__nor2_2
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08717_ _08718_/A _08718_/B vssd1 vssd1 vccd1 vccd1 _08717_/X sky130_fd_sc_hd__and2_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09693_/A _09690_/Y _09692_/B vssd1 vssd1 vccd1 vccd1 _09698_/B sky130_fd_sc_hd__o21ai_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08648_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _08649_/B sky130_fd_sc_hd__xnor2_1
XFILLER_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08555_/B _08579_/B vssd1 vssd1 vccd1 vccd1 _08579_/X sky130_fd_sc_hd__and2b_1
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _14997_/D sky130_fd_sc_hd__nor2_1
X_11590_ _11678_/A _11658_/A vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__nand2_1
XFILLER_179_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ _10609_/A _10541_/B vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__nand2_1
XFILLER_210_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _13259_/A _13297_/A _13259_/C vssd1 vssd1 vccd1 vccd1 _13261_/B sky130_fd_sc_hd__o21ai_1
XFILLER_41_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10472_ _10472_/A vssd1 vssd1 vccd1 vccd1 _14898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A _15475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ _12211_/A _12211_/B vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__xor2_1
XFILLER_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13191_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13195_/A sky130_fd_sc_hd__xnor2_1
XFILLER_151_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__A0 _15378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12142_ _12207_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__and2_1
XFILLER_68_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12073_ _12073_/A _12073_/B vssd1 vssd1 vccd1 vccd1 _12074_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11024_ _14923_/Q _14989_/Q vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10701__A _10701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08378__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15763_/CLK _15763_/D _14841_/Y vssd1 vssd1 vccd1 vccd1 _15763_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12976_/A _12976_/B _12976_/C vssd1 vssd1 vccd1 vccd1 _13690_/A sky130_fd_sc_hd__a21oi_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14714_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11926_ _11984_/B _11926_/B vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__xnor2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15694_ _15694_/CLK _15694_/D _14769_/Y vssd1 vssd1 vccd1 vccd1 _15694_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14645_/Y sky130_fd_sc_hd__inv_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11859_/C sky130_fd_sc_hd__xnor2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10808_ _15119_/Q _10103_/Y _10809_/C vssd1 vssd1 vccd1 vccd1 _14905_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14576_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14576_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11788_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__or2_1
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13527_ _13527_/A _13590_/A vssd1 vssd1 vccd1 vccd1 _15642_/D sky130_fd_sc_hd__xor2_1
X_10739_ _15714_/Q _15780_/Q vssd1 vssd1 vccd1 vccd1 _10741_/A sky130_fd_sc_hd__or2_1
XANTENNA__14843__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12066__C _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13458_ _13491_/S _13432_/B _13378_/B vssd1 vssd1 vccd1 vccd1 _13459_/B sky130_fd_sc_hd__o21a_1
XFILLER_51_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12409_ _12410_/A _12410_/C _12590_/A vssd1 vssd1 vccd1 vccd1 _12423_/A sky130_fd_sc_hd__o21a_1
XANTENNA_repeater701_A _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13389_ _13390_/A _13390_/B vssd1 vssd1 vccd1 vccd1 _13441_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ _15694_/CLK _15128_/D _14170_/Y vssd1 vssd1 vccd1 vccd1 _15128_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13178__B _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07950_ _15119_/Q _15284_/Q vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__nand2_1
X_15059_ _15107_/CLK _15059_/D _14097_/Y vssd1 vssd1 vccd1 vccd1 _15059_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07881_ _07881_/A vssd1 vssd1 vccd1 vccd1 _15327_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11707__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ _09778_/A _09551_/B vssd1 vssd1 vccd1 vccd1 _15171_/D sky130_fd_sc_hd__xor2_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08502_ _08500_/Y _08559_/B _12662_/A vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13922__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09482_ _09482_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _15280_/D sky130_fd_sc_hd__nor2_2
XFILLER_91_580 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ _08728_/B _08433_/B vssd1 vssd1 vccd1 vccd1 _08669_/A sky130_fd_sc_hd__xnor2_1
XFILLER_211_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08735__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08364_ _15041_/Q vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__buf_6
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ _11435_/A _11467_/A _08292_/B _08290_/B vssd1 vssd1 vccd1 vccd1 _08295_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14753__A _14753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15734__D _15734_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11617__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _09818_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _15744_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08198__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _15066_/Q _15099_/Q vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__and2b_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_912 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12760_ _12688_/A _12688_/B _12759_/X vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__a21boi_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A x_i_7[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11862_/A vssd1 vssd1 vccd1 vccd1 _11714_/A sky130_fd_sc_hd__inv_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A _13057_/A vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__or2b_2
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08645__B _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A _11352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14430_ _14435_/A vssd1 vssd1 vccd1 vccd1 _14430_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11642_ _11642_/A _11642_/B _11642_/C vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__nand3_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14361_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14361_/Y sky130_fd_sc_hd__inv_2
X_11573_ _11866_/A _11866_/B _11865_/C vssd1 vssd1 vccd1 vccd1 _12369_/C sky130_fd_sc_hd__a21o_1
XFILLER_126_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14663__A _14675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 x_i_0[9] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13312_ _13357_/B _13312_/B vssd1 vssd1 vccd1 vccd1 _13313_/B sky130_fd_sc_hd__or2_1
XANTENNA_input80_A x_i_4[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 x_i_1[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10524_ _10600_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _15026_/D sky130_fd_sc_hd__xor2_1
XFILLER_196_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14292_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14292_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ _13319_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13244_/C sky130_fd_sc_hd__xnor2_1
X_10455_ _10455_/A _10455_/B vssd1 vssd1 vccd1 vccd1 _14894_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08380__B _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13174_ _13247_/B _13216_/B vssd1 vssd1 vccd1 vccd1 _13722_/A sky130_fd_sc_hd__nand2_4
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10386_ _15104_/Q vssd1 vssd1 vccd1 vccd1 _10386_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12125_ _12183_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12128_/A sky130_fd_sc_hd__xnor2_4
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _12056_/A _12056_/B _12056_/C vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__and3_1
Xrepeater608 _11264_/X vssd1 vssd1 vccd1 vccd1 output476/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output334_A output334/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12630__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater619 repeater620/X vssd1 vssd1 vccd1 vccd1 output272/A sky130_fd_sc_hd__buf_4
X_11007_ _15278_/Q _11006_/Y _11005_/B vssd1 vssd1 vccd1 vccd1 _11008_/B sky130_fd_sc_hd__a21o_1
XFILLER_120_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15815_ _15815_/A vssd1 vssd1 vccd1 vccd1 _15815_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11246__B _15036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14838__A _14841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15746_ _15749_/CLK _15746_/D _14824_/Y vssd1 vssd1 vccd1 vccd1 _15746_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _13030_/C _13037_/B _13145_/A vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_794 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ _12254_/A _12247_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__nand2_1
XFILLER_179_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15677_ _15677_/CLK _15677_/D _14751_/Y vssd1 vssd1 vccd1 vccd1 _15677_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater651_A repeater653/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ _13357_/B _13201_/A _12888_/C vssd1 vssd1 vccd1 vccd1 _12923_/B sky130_fd_sc_hd__a21oi_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater749_A _15653_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14628_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14628_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14559_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14573__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater916_A input196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07886__S _07892_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _08290_/B _08087_/B _08088_/A _08079_/Y vssd1 vssd1 vccd1 vccd1 _08083_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08571__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__A _12451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__B _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__A1 _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13917__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A2 _15452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08982_ _15365_/Q _08983_/B _13591_/B vssd1 vssd1 vccd1 vccd1 _08986_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _15053_/Q _15218_/Q vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__nand2_1
XFILLER_190_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07864_ _15335_/Q _07864_/A1 _07900_/S vssd1 vssd1 vccd1 vccd1 _07865_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _09603_/A _09611_/A vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07795_ _15369_/Q _07795_/A1 _07795_/S vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10687__A_N _15279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14748__A _14750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _15539_/Q _15523_/Q _09533_/X vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _09465_/A _09473_/A vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nand2_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ _15043_/Q vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__buf_6
XFILLER_196_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09396_ _15410_/Q _15394_/Q vssd1 vssd1 vccd1 vccd1 _09398_/A sky130_fd_sc_hd__or2b_1
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08347_ _08347_/A _08347_/B _08347_/C vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__and3_1
XANTENNA__14483__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08278_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08314_/B sky130_fd_sc_hd__xnor2_1
XFILLER_192_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08481__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15729__D _15729_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10240_ _10239_/A _10239_/C _11406_/A vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__a21oi_1
XFILLER_191_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _10171_/A vssd1 vssd1 vccd1 vccd1 _15805_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08944__A2 _15448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput480 _11280_/X vssd1 vssd1 vccd1 vccd1 y_r_4[9] sky130_fd_sc_hd__buf_2
XFILLER_117_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput491 _15613_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[3] sky130_fd_sc_hd__buf_2
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10555__B_N _15295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ _13937_/A vssd1 vssd1 vccd1 vccd1 _13930_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input232_A x_r_6[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _13859_/A _13859_/B _13860_/A vssd1 vssd1 vccd1 vccd1 _13863_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14658__A _14660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15600_ _15768_/CLK _15600_/D _14670_/Y vssd1 vssd1 vccd1 vccd1 _15600_/Q sky130_fd_sc_hd__dfrtp_1
X_12812_ _12812_/A _12721_/B vssd1 vssd1 vccd1 vccd1 _12832_/B sky130_fd_sc_hd__or2b_1
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13792_ _13782_/B _13792_/B vssd1 vssd1 vccd1 vccd1 _13792_/X sky130_fd_sc_hd__and2b_1
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15531_ _15553_/CLK _15531_/D _14596_/Y vssd1 vssd1 vccd1 vccd1 _15531_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _13431_/B _12743_/B vssd1 vssd1 vccd1 vccd1 _12795_/A sky130_fd_sc_hd__nand2_1
XFILLER_128_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15493_/CLK _15462_/D _14524_/Y vssd1 vssd1 vccd1 vccd1 _15462_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11513__C _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _13145_/A _12970_/A vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__nand2_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14413_/Y sky130_fd_sc_hd__inv_2
X_11625_ _11624_/Y _11468_/B _11832_/A vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15393_ _15588_/CLK _15393_/D _14451_/Y vssd1 vssd1 vccd1 vccd1 _15393_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14393__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_85_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14344_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14344_/Y sky130_fd_sc_hd__inv_2
X_11556_ _12244_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_output284_A output284/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ _15255_/Q _15288_/Q vssd1 vssd1 vccd1 vccd1 _10508_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14275_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14275_/Y sky130_fd_sc_hd__inv_2
X_11487_ _11563_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__xnor2_1
XFILLER_183_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _13227_/B _13381_/B _13319_/A vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__and3_1
X_10438_ _10437_/A _10437_/C _10437_/B vssd1 vssd1 vccd1 vccd1 _10439_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_output451_A output451/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13157_ _13157_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__xnor2_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10369_ _10368_/A _10368_/B _10482_/A vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__a21oi_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__A _15051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12108_ _12308_/S _12108_/B vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__nand2_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13088_ _13089_/A _13089_/B vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__or2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater699_A _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _12110_/S _12178_/A _11959_/A _12038_/X vssd1 vssd1 vccd1 vccd1 _12040_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_867 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14568__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_53_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07580_ _07580_/A vssd1 vssd1 vccd1 vccd1 _15475_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_714 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15729_ _15729_/CLK _15729_/D _14806_/Y vssd1 vssd1 vccd1 vccd1 _15729_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12088__A _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09250_ _09250_/A _09250_/B _09250_/C vssd1 vssd1 vccd1 vccd1 _09250_/X sky130_fd_sc_hd__and3_1
XFILLER_178_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__xnor2_1
XFILLER_194_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09181_ _09188_/A _09189_/A vssd1 vssd1 vccd1 vccd1 _09654_/A sky130_fd_sc_hd__or2_1
XFILLER_147_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12816__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _11617_/A _11467_/A vssd1 vssd1 vccd1 vccd1 _08223_/C sky130_fd_sc_hd__xor2_1
XFILLER_175_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08063_ _08290_/B _08069_/B _08070_/B _08062_/X vssd1 vssd1 vccd1 vccd1 _08066_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput208 x_r_4[7] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__clkbuf_2
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _15196_/D sky130_fd_sc_hd__nor2_1
Xinput219 x_r_5[2] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07916_ _15525_/Q _15509_/Q vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__nand2_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08896_ _15470_/Q _15454_/Q vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__or2b_1
XFILLER_56_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater950 input148/X vssd1 vssd1 vccd1 vccd1 _07750_/A1 sky130_fd_sc_hd__buf_4
XFILLER_186_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1095 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater961 input133/X vssd1 vssd1 vccd1 vccd1 _07878_/A1 sky130_fd_sc_hd__clkbuf_2
X_07847_ _07847_/A vssd1 vssd1 vccd1 vccd1 _15344_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater972 repeater973/X vssd1 vssd1 vccd1 vccd1 _07388_/A1 sky130_fd_sc_hd__buf_4
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14478__A _14480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater983 input110/X vssd1 vssd1 vccd1 vccd1 _07532_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_204_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07778_ _07778_/A vssd1 vssd1 vccd1 vccd1 _15378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07380__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _09449_/A _09517_/B vssd1 vssd1 vccd1 vccd1 _09518_/C sky130_fd_sc_hd__and2b_1
XFILLER_17_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09448_ _15534_/Q _15518_/Q vssd1 vssd1 vccd1 vccd1 _09518_/A sky130_fd_sc_hd__and2_1
XFILLER_197_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09379_/A _09382_/B vssd1 vssd1 vccd1 vccd1 _09380_/A sky130_fd_sc_hd__and2_1
XFILLER_33_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11410_ _11411_/A _11411_/C _11411_/B vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12390_ _12390_/A _11728_/A vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__or2b_1
XFILLER_149_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ _11341_/A _11341_/B vssd1 vssd1 vccd1 vccd1 _11341_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input182_A x_r_3[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14060_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14060_/Y sky130_fd_sc_hd__inv_2
X_11272_ _11273_/A _11273_/B vssd1 vssd1 vccd1 vccd1 _11272_/X sky130_fd_sc_hd__xor2_4
XFILLER_165_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _13012_/A _13012_/B vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__nand2_1
X_10223_ _10221_/Y _10223_/B vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input43_A x_i_2[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _10155_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _15803_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14962_ _15694_/CLK _14962_/D _13994_/Y vssd1 vssd1 vccd1 vccd1 _14962_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10085_ _15116_/Q _15215_/Q vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__and2b_1
X_13913_ _15347_/Q _15331_/Q _13912_/X vssd1 vssd1 vccd1 vccd1 _13914_/B sky130_fd_sc_hd__a21o_1
X_14893_ _15792_/CLK _14893_/D _13922_/Y vssd1 vssd1 vccd1 vccd1 _14893_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14388__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ _13844_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13845_/A sky130_fd_sc_hd__and2_1
XFILLER_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08386__A _08396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13775_ _13775_/A _13862_/B vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__xnor2_2
X_10987_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _15011_/D sky130_fd_sc_hd__xor2_1
XFILLER_167_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15514_ _15749_/CLK _15514_/D _14578_/Y vssd1 vssd1 vccd1 vccd1 _15514_/Q sky130_fd_sc_hd__dfrtp_4
X_12726_ _12726_/A _12726_/B _12726_/C vssd1 vssd1 vccd1 vccd1 _12726_/X sky130_fd_sc_hd__or3_1
XFILLER_15_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output499_A _11212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15445_ _15558_/CLK _15445_/D _14506_/Y vssd1 vssd1 vccd1 vccd1 _15445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12657_ _12657_/A _12657_/B vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__or2_2
XFILLER_169_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__xor2_1
XFILLER_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15376_ _15617_/CLK _15376_/D _14432_/Y vssd1 vssd1 vccd1 vccd1 _15376_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08605__A1 _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _12588_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _15681_/D sky130_fd_sc_hd__xnor2_2
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08605__B2 _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14327_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14327_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11539_ _08123_/A _08123_/B _11462_/B _11432_/X vssd1 vssd1 vccd1 vccd1 _11828_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14851__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater614_A _10748_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14258_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14258_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _13722_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__xnor2_4
XFILLER_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14189_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14189_/Y sky130_fd_sc_hd__inv_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07701_ _07701_/A vssd1 vssd1 vccd1 vccd1 _15416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08681_ _13438_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14298__A _14299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A _11728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _15449_/Q _07632_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07563_ _15483_/Q _07563_/A1 _07579_/S vssd1 vssd1 vccd1 vccd1 _07564_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09302_ _15404_/Q _15388_/Q vssd1 vssd1 vccd1 vccd1 _09302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13930__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _15517_/Q _07494_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _09233_/A _09233_/B vssd1 vssd1 vccd1 vccd1 _15239_/D sky130_fd_sc_hd__xor2_2
XFILLER_181_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09164_ _15565_/Q _15545_/Q _09160_/B vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__o21a_1
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _08120_/C _08115_/B vssd1 vssd1 vccd1 vccd1 _08325_/B sky130_fd_sc_hd__xnor2_2
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ _15500_/Q _15484_/Q vssd1 vssd1 vccd1 vccd1 _09095_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14761__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_731 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08046_ _08064_/A _08064_/B _08045_/Y vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13353__B1 _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14911__D _14911_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_680 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_627 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _09997_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _14933_/D sky130_fd_sc_hd__xor2_1
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07583__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _15466_/Q _15450_/Q _08947_/B vssd1 vssd1 vccd1 vccd1 _08948_/X sky130_fd_sc_hd__o21a_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A2 _15391_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13824__B _13824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08879_ _15467_/Q _15451_/Q vssd1 vssd1 vccd1 vccd1 _08879_/X sky130_fd_sc_hd__and2b_1
XANTENNA__15742__D _15742_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10910_ _10910_/A _11119_/A _10910_/C vssd1 vssd1 vccd1 vccd1 _10912_/A sky130_fd_sc_hd__and3_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater780 repeater781/X vssd1 vssd1 vccd1 vccd1 output494/A sky130_fd_sc_hd__buf_4
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater791 repeater792/X vssd1 vssd1 vccd1 vccd1 output461/A sky130_fd_sc_hd__buf_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _11890_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__nand2_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14001__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ _10839_/X _10843_/C vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__and2b_1
XFILLER_60_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13560_ _13560_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13561_/C sky130_fd_sc_hd__or2_1
X_10772_ _15720_/Q _15786_/Q vssd1 vssd1 vccd1 vccd1 _11287_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12631__A2 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12511_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13491_ _13432_/B _13432_/A _13491_/S vssd1 vssd1 vccd1 vccd1 _13492_/B sky130_fd_sc_hd__mux2_2
XANTENNA__08653__B _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _15506_/CLK _15230_/D _14278_/Y vssd1 vssd1 vccd1 vccd1 _15230_/Q sky130_fd_sc_hd__dfrtp_1
X_12442_ _14947_/Q vssd1 vssd1 vccd1 vccd1 _12444_/A sky130_fd_sc_hd__inv_2
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15161_ _15180_/CLK _15161_/D _14205_/Y vssd1 vssd1 vccd1 vccd1 _15161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_614 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12373_ _12373_/A _12381_/B _12381_/C vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__and3_1
XANTENNA__14671__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14112_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14112_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11324_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11324_/X sky130_fd_sc_hd__xor2_2
XFILLER_158_1035 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15092_ _15110_/CLK _15092_/D _14132_/Y vssd1 vssd1 vccd1 vccd1 _15092_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14043_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14043_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11255_ _15711_/Q _11254_/Y _11253_/B vssd1 vssd1 vccd1 vccd1 _11257_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12191__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_73 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10206_ _11396_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11186_/A _11186_/B vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__nand2_4
XFILLER_45_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11370__A2 _15029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ _10135_/Y _10137_/B vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__nand2b_2
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14945_ _15791_/CLK _14945_/D _13976_/Y vssd1 vssd1 vccd1 vccd1 _14945_/Q sky130_fd_sc_hd__dfrtp_1
X_10068_ _15213_/Q _15114_/Q vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__and2b_1
XANTENNA_output414_A output414/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15652__D _15652_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14876_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13827_ _14976_/Q _13827_/B vssd1 vssd1 vccd1 vccd1 _13827_/X sky130_fd_sc_hd__and2_1
XANTENNA_repeater564_A repeater565/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14846__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13758_ _13754_/Y _13757_/X _13752_/B vssd1 vssd1 vccd1 vccd1 _13758_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ _12921_/A _12630_/A _12708_/X vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__a21o_1
XFILLER_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater731_A _15676_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13689_ _13700_/A _13700_/B vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_repeater829_A repeater830/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15428_ _15428_/CLK _15428_/D _14488_/Y vssd1 vssd1 vccd1 vccd1 _15428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_1050 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _15717_/CLK _15359_/D _14414_/Y vssd1 vssd1 vccd1 vccd1 _15359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07894__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13909__B _15330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _14962_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07907__B _15445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13886__A1 _15338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_907 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _09851_/A vssd1 vssd1 vccd1 vccd1 _15752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A1 _07565_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08802_ _08802_/A vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13925__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09552_/Y _09781_/B _09554_/B vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__o21ai_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08733_ _12810_/A _12780_/A _08731_/X _08732_/Y vssd1 vssd1 vccd1 vccd1 _08733_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11445__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08664_ _12703_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__and2_1
XFILLER_96_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _07615_/A vssd1 vssd1 vccd1 vccd1 _15458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08598_/A _08621_/A vssd1 vssd1 vccd1 vccd1 _08596_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14756__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ _07546_/A vssd1 vssd1 vccd1 vccd1 _15492_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08754__A _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09569__B _15419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ _15525_/Q _07477_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09216_ _09211_/A _09215_/B _09211_/B vssd1 vssd1 vccd1 vccd1 _15300_/D sky130_fd_sc_hd__o21ba_1
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ _09147_/A _09147_/B vssd1 vssd1 vccd1 vccd1 _15285_/D sky130_fd_sc_hd__nor2_1
XANTENNA__14491__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _15496_/Q _15480_/Q vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15737__D _15737_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08029_ _11458_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08097_/B sky130_fd_sc_hd__xor2_2
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11040_ _11032_/Y _11036_/B _11034_/B vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__o21ai_1
XFILLER_157_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input145_A x_r_0[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08929__A _15476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A _12991_/B vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__or2_1
XFILLER_188_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _14739_/A vssd1 vssd1 vccd1 vccd1 _14730_/Y sky130_fd_sc_hd__inv_2
X_11942_ _15733_/Q _11950_/B vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14661_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _12544_/A _11873_/B vssd1 vssd1 vccd1 vccd1 _11945_/B sky130_fd_sc_hd__and2b_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14666__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13612_/A _13613_/B vssd1 vssd1 vccd1 vccd1 _15095_/D sky130_fd_sc_hd__xnor2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12065__B1 _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10824_ _10823_/B _10823_/C _10823_/A vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__a21oi_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14592_/Y sky130_fd_sc_hd__inv_2
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _13543_/A _13546_/B vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__and2_1
XFILLER_201_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10755_ _15717_/Q _15783_/Q vssd1 vssd1 vccd1 vccd1 _10756_/B sky130_fd_sc_hd__nand2_1
XFILLER_203_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__A2 _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ _13781_/A _13781_/B vssd1 vssd1 vccd1 vccd1 _13771_/B sky130_fd_sc_hd__xor2_4
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10686_ _15278_/Q _15179_/Q vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15213_ _15460_/CLK _15213_/D _14261_/Y vssd1 vssd1 vccd1 vccd1 _15213_/Q sky130_fd_sc_hd__dfrtp_1
X_12425_ _14945_/Q _12425_/B vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__and2_1
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12914__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ _15394_/CLK _15144_/D _14187_/Y vssd1 vssd1 vccd1 vccd1 _15144_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12356_ _12358_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__xnor2_4
XFILLER_5_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput309 output309/A vssd1 vssd1 vccd1 vccd1 y_i_2[8] sky130_fd_sc_hd__buf_2
XANTENNA_output364_A output364/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07795__A1 _07795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _14923_/Q _11306_/Y _11305_/B vssd1 vssd1 vccd1 vccd1 _11309_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15075_ _15750_/CLK _15075_/D _14114_/Y vssd1 vssd1 vccd1 vccd1 _15075_/Q sky130_fd_sc_hd__dfrtp_1
X_12287_ _12287_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__nor2_1
X_14026_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14026_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11238_ _15034_/Q vssd1 vssd1 vccd1 vccd1 _11238_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output531_A _15635_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _11169_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11169_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08839__A _15348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_556 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater681_A _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater779_A _15618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13183__C _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ _15192_/CLK _14928_/D _13959_/Y vssd1 vssd1 vccd1 vccd1 _14928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_656 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14859_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14859_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater946_A input152/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_998 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14576__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ _15567_/Q _07400_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08380_ _12945_/A _12881_/A vssd1 vssd1 vccd1 vccd1 _08422_/C sky130_fd_sc_hd__xor2_1
XFILLER_1_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_470 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_694 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _13600_/A _08998_/B _09000_/X vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__a21o_1
XFILLER_178_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15557__D input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_734 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09903_ _15223_/Q _15190_/Q vssd1 vssd1 vccd1 vccd1 _09904_/C sky130_fd_sc_hd__or2b_1
XFILLER_63_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07538__A1 input107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09834_ _09834_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _15748_/D sky130_fd_sc_hd__nor2_2
XFILLER_63_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ _15101_/Q _15068_/Q vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__and2b_1
XFILLER_6_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08716_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08718_/A sky130_fd_sc_hd__inv_2
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_399 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09696_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__nand2_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _12810_/A _08369_/B _08646_/Y vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__a21oi_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14486__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__A1 input216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13390__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07799__S _07803_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08577_/A _08564_/Y _08631_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08586_/B
+ sky130_fd_sc_hd__o22ai_4
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11622__B _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ _07529_/A vssd1 vssd1 vccd1 vccd1 _15500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10540_ _15260_/Q _15293_/Q vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10469_/X _10473_/C vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__and2b_1
XFILLER_41_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _12149_/A _12150_/A _12149_/B _12209_/X vssd1 vssd1 vccd1 vccd1 _12211_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_157_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13190_ _13263_/A _13190_/B vssd1 vssd1 vccd1 vccd1 _13249_/B sky130_fd_sc_hd__or2_1
XFILLER_68_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07777__A1 _07777_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12141_ _12141_/A _12141_/B _12141_/C vssd1 vssd1 vccd1 vccd1 _12142_/B sky130_fd_sc_hd__or3_1
XFILLER_124_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12072_ _12132_/S _12204_/A _11990_/A _12071_/X vssd1 vssd1 vccd1 vccd1 _12073_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ _14923_/Q _14989_/Q vssd1 vssd1 vccd1 vccd1 _11023_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08378__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _13052_/B _12974_/B vssd1 vssd1 vccd1 vccd1 _12976_/C sky130_fd_sc_hd__xor2_4
X_15762_ _15763_/CLK _15762_/D _14840_/Y vssd1 vssd1 vccd1 vccd1 _15762_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14713_/Y sky130_fd_sc_hd__inv_2
X_11925_ _11835_/A _11835_/B _11848_/B _11853_/A vssd1 vssd1 vccd1 vccd1 _11926_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15693_/CLK _15693_/D _14768_/Y vssd1 vssd1 vccd1 vccd1 _15693_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14396__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _11931_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__and2_1
XFILLER_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14644_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14644_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08394__A _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__S _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_930 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10807_ _10104_/Y _15284_/Q _10103_/B vssd1 vssd1 vccd1 vccd1 _10809_/C sky130_fd_sc_hd__a21o_1
X_14575_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14575_/Y sky130_fd_sc_hd__inv_2
X_11787_ _15731_/Q _11787_/B _11787_/C vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__and3_1
XANTENNA__13808__B_N _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10738_ _11259_/A _10738_/B vssd1 vssd1 vccd1 vccd1 _10738_/Y sky130_fd_sc_hd__xnor2_1
X_13526_ _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__xnor2_2
XFILLER_207_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13457_ _13433_/Y _13432_/A _13456_/Y vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__a21oi_1
XFILLER_51_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10669_ _10990_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_173_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _14944_/Q _12591_/B vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__xnor2_2
XFILLER_127_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _13386_/X _13441_/A vssd1 vssd1 vccd1 vccd1 _13390_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15127_ _15433_/CLK _15127_/D _14169_/Y vssd1 vssd1 vccd1 vccd1 _15127_/Q sky130_fd_sc_hd__dfrtp_1
X_12339_ _15741_/Q _12339_/B vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__or2_1
XFILLER_154_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ _15107_/CLK _15058_/D _14096_/Y vssd1 vssd1 vccd1 vccd1 _15058_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater896_A input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14009_/Y sky130_fd_sc_hd__inv_2
X_07880_ _15327_/Q input132/X _07892_/S vssd1 vssd1 vccd1 vccd1 _07881_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08569__A _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10611__B _15294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ _09549_/Y _15415_/Q _09547_/B vssd1 vssd1 vccd1 vccd1 _09551_/B sky130_fd_sc_hd__a21o_1
XFILLER_209_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08501_ _15792_/Q _12688_/A vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__xor2_2
XFILLER_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ _09480_/A _09480_/B _09529_/A vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__a21oi_1
XFILLER_184_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ _08432_/A _08666_/A vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__xnor2_1
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07412__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08363_ _12881_/A _12654_/A vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ _11707_/A vssd1 vssd1 vccd1 vccd1 _11545_/A sky130_fd_sc_hd__inv_2
XFILLER_108_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07759__A1 _07759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10074__A _10074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08479__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09817_ _09816_/A _09816_/C _09816_/B vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__a21oi_1
XFILLER_86_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08198__B _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09748_ _15065_/Q _15098_/Q vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__nand2_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09678_/Y _15555_/Q _09677_/B vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_924 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11710_ _11710_/A _11710_/B vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__or2_1
XFILLER_14_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12690_/A _12690_/B _12690_/C vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__nand3_1
XANTENNA_input108_A x_i_6[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11641_ _11642_/A _11642_/B _11642_/C vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__a21oi_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14360_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__buf_8
XFILLER_211_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _11866_/A _11865_/C _11866_/B vssd1 vssd1 vccd1 vccd1 _12369_/B sky130_fd_sc_hd__nand3_1
XFILLER_195_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13311_ _13357_/B _13312_/B vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 x_i_1[0] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
X_10523_ _10598_/A _10518_/B _10522_/X vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__a21o_1
XFILLER_183_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14291_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ _13240_/X _13340_/A vssd1 vssd1 vccd1 vccd1 _13319_/B sky130_fd_sc_hd__and2b_1
XFILLER_182_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10454_ _10453_/B _10453_/C _10453_/A vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_input73_A x_i_4[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ _13173_/A _13173_/B _13173_/C vssd1 vssd1 vccd1 vccd1 _13216_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10385_ _10385_/A _10385_/B vssd1 vssd1 vccd1 vccd1 _14940_/D sky130_fd_sc_hd__nor2_1
XFILLER_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12124_ _12055_/A _12055_/B _12054_/A vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__13295__A _13737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12056_/C sky130_fd_sc_hd__xnor2_1
XFILLER_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater609 _11175_/X vssd1 vssd1 vccd1 vccd1 output510/A sky130_fd_sc_hd__clkbuf_2
X_11006_ _15179_/Q vssd1 vssd1 vccd1 vccd1 _11006_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12630__C _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output327_A _15669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ _15814_/A vssd1 vssd1 vccd1 vccd1 _15814_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15745_ _15749_/CLK _15745_/D _14823_/Y vssd1 vssd1 vccd1 vccd1 _15745_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A _12970_/A _13046_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__and3_1
XANTENNA__15660__D _15660_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12639__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__nand2_1
XFILLER_179_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15676_ _15707_/CLK _15676_/D _14750_/Y vssd1 vssd1 vccd1 vccd1 _15676_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _13357_/B _13201_/A _12888_/C vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__and3_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09013__A _15373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14627_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14627_/Y sky130_fd_sc_hd__inv_2
X_11839_ _12254_/A _12144_/A _11839_/C vssd1 vssd1 vccd1 vccd1 _12002_/B sky130_fd_sc_hd__and3_1
XANTENNA_repeater644_A _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14854__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14558_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14558_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08852__A _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13803_/A _13519_/B vssd1 vssd1 vccd1 vccd1 _13791_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_repeater811_A repeater812/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14489_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08571__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ _08986_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _13591_/B sky130_fd_sc_hd__or2_1
XFILLER_103_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11718__A _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ _07932_/A vssd1 vssd1 vccd1 vccd1 _14921_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07915__B _15381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07863_ _07863_/A vssd1 vssd1 vccd1 vccd1 _15336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _15441_/Q _15425_/Q vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13933__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ _07794_/A vssd1 vssd1 vccd1 vccd1 _15370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08879__A_N _15467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09533_ _15539_/Q _15523_/Q _09532_/B vssd1 vssd1 vccd1 vccd1 _09533_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09464_ _15536_/Q _15520_/Q vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__or2b_1
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _12945_/A _12881_/A vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__nand2_1
X_09395_ _09397_/A _09397_/B vssd1 vssd1 vccd1 vccd1 _15148_/D sky130_fd_sc_hd__xor2_1
XANTENNA__14764__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08346_ _08322_/A _08322_/B _08324_/Y _08345_/Y vssd1 vssd1 vccd1 vccd1 _08347_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _08277_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08277_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_164_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10170_ _10168_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__and2b_1
XFILLER_65_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13827__B _13827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput470 output470/A vssd1 vssd1 vccd1 vccd1 y_r_4[15] sky130_fd_sc_hd__buf_2
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15745__D _15745_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput481 _15815_/X vssd1 vssd1 vccd1 vccd1 y_r_5[0] sky130_fd_sc_hd__buf_2
XANTENNA__11628__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput492 _15614_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[4] sky130_fd_sc_hd__buf_2
XANTENNA__14004__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08002__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _13860_/A _13860_/B vssd1 vssd1 vccd1 vccd1 _15673_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_input225_A x_r_5[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08897__B_N _15471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A _15462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _12811_/A _12811_/B vssd1 vssd1 vccd1 vccd1 _12832_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _13791_/A _13791_/B vssd1 vssd1 vccd1 vccd1 _13794_/A sky130_fd_sc_hd__xnor2_1
XFILLER_15_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15530_ _15542_/CLK _15530_/D _14595_/Y vssd1 vssd1 vccd1 vccd1 _15530_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12781_/A _12781_/B vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__xor2_1
XFILLER_63_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _14919_/Q vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__clkbuf_4
X_15461_ _15700_/CLK _15461_/D _14523_/Y vssd1 vssd1 vccd1 vccd1 _15461_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_179_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11624_ _11906_/A vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__clkinv_2
X_14412_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14412_/Y sky130_fd_sc_hd__inv_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15392_ _15392_/CLK _15392_/D _14450_/Y vssd1 vssd1 vccd1 vccd1 _15392_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08672__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12964__A1 _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ _11555_/A _11623_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__xnor2_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14343_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14343_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ _15255_/Q _15288_/Q vssd1 vssd1 vccd1 vccd1 _10506_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14274_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14274_/Y sky130_fd_sc_hd__inv_2
X_11486_ _11564_/A _11564_/B vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output277_A output277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13225_ _13320_/A _13321_/A vssd1 vssd1 vccd1 vccd1 _13231_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12932__A1_N _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10437_ _10437_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__and3_1
XFILLER_124_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156_ _13235_/B _13156_/B vssd1 vssd1 vccd1 vccd1 _13157_/B sky130_fd_sc_hd__xnor2_1
XFILLER_174_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10368_ _10368_/A _10368_/B _10482_/A vssd1 vssd1 vccd1 vccd1 _10370_/A sky130_fd_sc_hd__and3_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13737__B _13737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output444_A output444/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ _12231_/A _12228_/A vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__nand2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13002_/A _13002_/B _13086_/Y vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__a21oi_1
X_10299_ _15121_/Q _15154_/Q vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12038_ _12038_/A _12038_/B vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__or2_1
XANTENNA__11257__B _11257_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater594_A _11367_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14849__A _14853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_879 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__A _15445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater761_A _15641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13989_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__A0 _15436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15728_ _15729_/CLK _15728_/D _14805_/Y vssd1 vssd1 vccd1 vccd1 _15728_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15659_ _15699_/CLK _15659_/D _14732_/Y vssd1 vssd1 vccd1 vccd1 _15659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14584__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08200_ _15014_/Q vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__buf_6
XFILLER_178_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ _15570_/Q _15550_/Q vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__and2_1
XFILLER_187_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12816__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _15006_/Q vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_175_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12308__S _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08062_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__or2_1
XFILLER_146_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13928__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput209 x_r_4[8] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_2
X_08964_ _08963_/B _08963_/C _08963_/A vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__o21a_1
XFILLER_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _15397_/Q _15381_/Q vssd1 vssd1 vccd1 vccd1 _15119_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08895_ _08957_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14759__A _14761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07898__A0 _15318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater940 repeater941/X vssd1 vssd1 vccd1 vccd1 _07757_/A1 sky130_fd_sc_hd__buf_6
X_07846_ _15344_/Q input197/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater951 input147/X vssd1 vssd1 vccd1 vccd1 _07771_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater962 input13/X vssd1 vssd1 vccd1 vccd1 _07632_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater973 input118/X vssd1 vssd1 vccd1 vccd1 repeater973/X sky130_fd_sc_hd__buf_2
XFILLER_186_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater984 input105/X vssd1 vssd1 vccd1 vccd1 _07512_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07777_ _15378_/Q _07777_/A1 _07791_/S vssd1 vssd1 vccd1 vccd1 _07778_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14909__D _14909_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08476__B _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ _09516_/A _09517_/B vssd1 vssd1 vccd1 vccd1 _15260_/D sky130_fd_sc_hd__xnor2_1
XFILLER_25_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _15534_/Q _15518_/Q vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__nor2_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14494__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ _09377_/B _09377_/C _09377_/A vssd1 vssd1 vccd1 vccd1 _09382_/B sky130_fd_sc_hd__o21ai_1
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07600__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08329_/X sky130_fd_sc_hd__and2_1
XFILLER_32_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07822__A0 _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _11339_/A _11339_/C _11339_/B vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _15715_/Q _11270_/Y _11269_/B vssd1 vssd1 vccd1 vccd1 _11273_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input175_A x_r_2[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ _13008_/X _13097_/A vssd1 vssd1 vccd1 vccd1 _13012_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10222_ _15075_/Q _15240_/Q vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13557__B _13563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ _15146_/Q _15311_/Q vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__xor2_2
XFILLER_82_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A x_i_2[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _15383_/CLK _14961_/D _13993_/Y vssd1 vssd1 vccd1 vccd1 _14961_/Q sky130_fd_sc_hd__dfrtp_1
X_10084_ _15215_/Q _15116_/Q vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__and2b_1
XFILLER_181_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14669__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13912_ _15347_/Q _15331_/Q _13911_/B vssd1 vssd1 vccd1 vccd1 _13912_/X sky130_fd_sc_hd__o21a_1
X_14892_ _15792_/CLK _14892_/D _13921_/Y vssd1 vssd1 vccd1 vccd1 _14892_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13843_ _13842_/B _13842_/C _13842_/A vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08386__B _12654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__A _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10986_ _15273_/Q _10985_/Y _10984_/B vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ _13774_/A _13774_/B vssd1 vssd1 vccd1 vccd1 _13862_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ _15542_/CLK _15513_/D _14577_/Y vssd1 vssd1 vccd1 vccd1 _15513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12725_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__xnor2_1
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15444_ _15444_/CLK _15444_/D _14505_/Y vssd1 vssd1 vccd1 vccd1 _15444_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ _12703_/A _12703_/B _12703_/C vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_output394_A output394/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07510__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11607_ _11607_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__xnor2_1
X_12587_ _12585_/A _12385_/B _12585_/B _12383_/Y vssd1 vssd1 vccd1 vccd1 _12588_/B
+ sky130_fd_sc_hd__a31o_1
X_15375_ _15375_/CLK _15375_/D _14431_/Y vssd1 vssd1 vccd1 vccd1 _15375_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14326_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14326_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ _11538_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11827_/C sky130_fd_sc_hd__nor2_1
XFILLER_184_784 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11469_ _11469_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11469_/Y sky130_fd_sc_hd__nand2_1
X_14257_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14257_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater607_A _11316_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _13208_/A _13208_/B vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__xnor2_4
X_14188_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14188_/Y sky130_fd_sc_hd__inv_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _13558_/B _15765_/Q vssd1 vssd1 vccd1 vccd1 _13213_/B sky130_fd_sc_hd__or2b_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14579__A _14580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater976_A input116/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _15416_/Q _07700_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08680_ _08680_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__xnor2_1
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07631_ _07631_/A vssd1 vssd1 vccd1 vccd1 _15450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07562_ _07562_/A vssd1 vssd1 vccd1 vccd1 _15484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09301_ _09368_/A _09301_/B vssd1 vssd1 vccd1 vccd1 _15125_/D sky130_fd_sc_hd__xnor2_1
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ _07493_/A vssd1 vssd1 vccd1 vccd1 _15518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09232_ _09230_/A _09230_/B _09231_/X vssd1 vssd1 vccd1 vccd1 _09233_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07420__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _09161_/Y _09163_/B vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__nand2b_1
X_08114_ _08112_/A _08112_/B _08120_/B vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__a21oi_1
XFILLER_147_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09094_ _09236_/A _09094_/B vssd1 vssd1 vccd1 vccd1 _15224_/D sky130_fd_sc_hd__xnor2_1
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _08045_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13353__A1 _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10082__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _15196_/Q _15229_/Q _09995_/B vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__a21o_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _08947_/A _08947_/B vssd1 vssd1 vccd1 vccd1 _15190_/D sky130_fd_sc_hd__xnor2_1
XFILLER_192_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14489__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11906__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08487__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _15468_/Q _15452_/Q vssd1 vssd1 vccd1 vccd1 _08952_/A sky130_fd_sc_hd__xnor2_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater770 _15628_/Q vssd1 vssd1 vccd1 vccd1 output524/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _07829_/A vssd1 vssd1 vccd1 vccd1 _15353_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater781 _15616_/Q vssd1 vssd1 vccd1 vccd1 repeater781/X sky130_fd_sc_hd__buf_2
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater792 _15601_/Q vssd1 vssd1 vccd1 vccd1 repeater792/X sky130_fd_sc_hd__buf_2
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _10839_/B _10839_/C _10839_/A vssd1 vssd1 vccd1 vccd1 _10843_/C sky130_fd_sc_hd__a21o_1
XFILLER_77_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_99_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _10768_/A _11283_/A _10768_/B _10770_/X vssd1 vssd1 vccd1 vccd1 _10774_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _14952_/Q _12510_/B vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nand2_1
X_13490_ _13490_/A _13490_/B vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__nor2_2
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ _12440_/A _12440_/C _12455_/C vssd1 vssd1 vccd1 vccd1 _12463_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__09111__A _15503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12372_/A _12372_/B vssd1 vssd1 vccd1 vccd1 _12381_/C sky130_fd_sc_hd__nand2_1
X_15160_ _15694_/CLK _15160_/D _14204_/Y vssd1 vssd1 vccd1 vccd1 _15160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14111_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14111_/Y sky130_fd_sc_hd__inv_2
X_11323_ _14927_/Q _11322_/Y _11321_/B vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__a21o_1
X_15091_ _15107_/CLK _15091_/D _14131_/Y vssd1 vssd1 vccd1 vccd1 _15091_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_180_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1047 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14042_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _15777_/Q vssd1 vssd1 vccd1 vccd1 _11254_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08161__S _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13287__B _13567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__B _15281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11088__A _11088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _11396_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _15761_/D sky130_fd_sc_hd__xor2_2
X_11185_ _15749_/Q _15027_/Q vssd1 vssd1 vccd1 vccd1 _11186_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _15143_/Q _15308_/Q vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14399__A _14399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14944_ _15791_/CLK _14944_/D _13975_/Y vssd1 vssd1 vccd1 vccd1 _14944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10067_ _15212_/Q _15113_/Q vssd1 vssd1 vccd1 vccd1 _10071_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14875_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14875_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output407_A output407/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ _13826_/A _13826_/B vssd1 vssd1 vccd1 vccd1 _13826_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ _13849_/B _13849_/C _14981_/Q vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_136_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15511_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10969_ _15170_/Q vssd1 vssd1 vccd1 vccd1 _10969_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11551__A _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ _12708_/A _12881_/A _12810_/A vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__and3_1
XFILLER_176_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13688_ _13688_/A _13688_/B _12976_/C vssd1 vssd1 vccd1 vccd1 _13700_/B sky130_fd_sc_hd__or3b_2
XFILLER_188_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15427_ _15428_/CLK _15427_/D _14487_/Y vssd1 vssd1 vccd1 vccd1 _15427_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_54_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12639_ _13012_/A _13201_/A vssd1 vssd1 vccd1 vccd1 _12813_/C sky130_fd_sc_hd__xor2_1
XANTENNA_repeater724_A repeater725/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14862__A _14862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1062 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09956__A _09956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _15364_/CLK _15358_/D _14413_/Y vssd1 vssd1 vccd1 vccd1 _15358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_795 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14309_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14309_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15289_ _15553_/CLK _15289_/D _14341_/Y vssd1 vssd1 vccd1 vccd1 _15289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13886__A2 _15322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _09848_/X _09852_/C vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__and2b_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08762__A1 _15333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08801_/A _13897_/A vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__or2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _15156_/D sky130_fd_sc_hd__xor2_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08732_ _08732_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _08732_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10630__A _15268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14102__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08663_ _08663_/A _08663_/B _08663_/C vssd1 vssd1 vccd1 vccd1 _08664_/B sky130_fd_sc_hd__or3_1
XFILLER_39_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13941__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ _15458_/Q input7/X _07632_/S vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__mux2_1
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__or2_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07545_ _15492_/Q _07545_/A1 _07589_/S vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_127_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07476_ _07476_/A vssd1 vssd1 vccd1 vccd1 _15526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _09680_/A _09215_/B vssd1 vssd1 vccd1 vccd1 _15299_/D sky130_fd_sc_hd__xor2_2
XFILLER_10_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14772__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09146_ _15561_/Q _15541_/Q _09628_/C vssd1 vssd1 vccd1 vccd1 _09147_/B sky130_fd_sc_hd__and3_1
XFILLER_33_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ _09077_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _15220_/D sky130_fd_sc_hd__xnor2_1
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08028_ _11458_/A vssd1 vssd1 vccd1 vccd1 _11447_/C sky130_fd_sc_hd__inv_2
XFILLER_123_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _09979_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _14926_/D sky130_fd_sc_hd__xnor2_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12841_/A _12987_/X _12989_/X _13690_/B vssd1 vssd1 vccd1 vccd1 _13290_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14012__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input138_A x_r_0[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _12455_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11950_/B sky130_fd_sc_hd__xnor2_2
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08010__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14660_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__inv_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11873_/B _12544_/A vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__and2b_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _09013_/Y _13610_/B _09015_/B vssd1 vssd1 vccd1 vccd1 _13613_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12065__A1 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _10823_/A _10823_/B _10823_/C vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__and3_1
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14591_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14591_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_118_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15249_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13542_ _13538_/Y _13536_/A _13536_/B _13539_/Y _13541_/A vssd1 vssd1 vccd1 vccd1
+ _13546_/B sky130_fd_sc_hd__a311o_1
XANTENNA__10615__A2 _15295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ _15717_/Q _15783_/Q vssd1 vssd1 vccd1 vccd1 _10754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__B _15001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07492__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10685_ _10685_/A _11003_/B vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__nand2_1
X_13473_ _13473_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13781_/B sky130_fd_sc_hd__xnor2_4
XFILLER_51_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15212_ _15460_/CLK _15212_/D _14259_/Y vssd1 vssd1 vccd1 vccd1 _15212_/Q sky130_fd_sc_hd__dfrtp_2
X_12424_ _12435_/A _12424_/B vssd1 vssd1 vccd1 vccd1 _15650_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ _15394_/CLK _15143_/D _14186_/Y vssd1 vssd1 vccd1 vccd1 _15143_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13298__A _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__xnor2_4
XFILLER_5_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ _14989_/Q vssd1 vssd1 vccd1 vccd1 _11306_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12286_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15074_ _15345_/CLK _15074_/D _14113_/Y vssd1 vssd1 vccd1 vccd1 _15074_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14025_/Y sky130_fd_sc_hd__inv_2
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11237_/Y sky130_fd_sc_hd__nor2_2
XFILLER_206_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11168_ _11167_/A _11167_/C _11359_/A vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output524_A output524/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15663__D _15663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08839__B _15332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _10817_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _15796_/D sky130_fd_sc_hd__xor2_1
XFILLER_132_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11350_/A sky130_fd_sc_hd__nor2_2
XFILLER_95_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ _15221_/CLK _14927_/D _13957_/Y vssd1 vssd1 vccd1 vccd1 _14927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14857__A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14858_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14858_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__xor2_4
XFILLER_91_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater841_A repeater842/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15773_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14789_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14789_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07483__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14592__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ _15369_/Q _15353_/Q vssd1 vssd1 vccd1 vccd1 _09000_/X sky130_fd_sc_hd__and2b_1
XFILLER_192_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_129_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09902_ _09900_/Y _09902_/B vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13936__A _13937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12840__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09833_ _09832_/B _09832_/C _09832_/A vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__a21oi_1
XFILLER_154_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09764_ _15068_/Q _15101_/Q vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__and2b_1
XFILLER_6_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08715_ _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _08715_/Y sky130_fd_sc_hd__nand2_1
X_09695_ _15056_/Q _15089_/Q vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14767__A _14774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ _12881_/A _12810_/A vssd1 vssd1 vccd1 vccd1 _08646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14917__D _14917_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__xor2_2
XFILLER_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11191__A _15750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07528_ _15500_/Q _07528_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07529_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11622__C _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07459_ _15534_/Q _07459_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _10469_/B _10469_/C _10469_/A vssd1 vssd1 vccd1 vccd1 _10473_/C sky130_fd_sc_hd__a21o_1
XANTENNA__15748__D _15748_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09129_/A _09265_/A vssd1 vssd1 vccd1 vccd1 _15231_/D sky130_fd_sc_hd__xor2_1
XFILLER_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14007__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12140_ _12141_/A _12141_/B _12141_/C vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08974__A1 _15475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08005__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12071_ _12071_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__or2_1
XANTENNA_input255_A x_r_7[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11022_ _14922_/Q _14988_/Q _11021_/Y _10861_/Y vssd1 vssd1 vccd1 vccd1 _11026_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_173_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15761_/CLK _15761_/D _14839_/Y vssd1 vssd1 vccd1 vccd1 _15761_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12973_ _12973_/A _12973_/B vssd1 vssd1 vccd1 vccd1 _12974_/B sky130_fd_sc_hd__nor2_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14677__A _14680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14712_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11924_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__xor2_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15692_ _15699_/CLK _15692_/D _14767_/Y vssd1 vssd1 vccd1 vccd1 _15692_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14643_ _14661_/A vssd1 vssd1 vccd1 vccd1 _14643_/Y sky130_fd_sc_hd__inv_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11855_/A _11855_/B _11855_/C vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__nand3_1
XFILLER_32_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_960 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _10806_/A _11300_/A vssd1 vssd1 vccd1 vccd1 _10806_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_198_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14574_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14574_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_942 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_621 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _15731_/Q _12541_/B vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__nor2_1
XFILLER_159_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13525_ _15774_/Q _13804_/B vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07465__A1 _07465_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ _10731_/A _10733_/B _10731_/B vssd1 vssd1 vccd1 vccd1 _10738_/B sky130_fd_sc_hd__a21boi_2
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12925__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A_N _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _13491_/S _13432_/B _13432_/A vssd1 vssd1 vccd1 vccd1 _13456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10668_ _10662_/A _10664_/B _10662_/B vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__a21boi_2
XANTENNA_output474_A _11256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ _12455_/D _12407_/B vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__or2_2
XFILLER_127_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10599_ _10515_/A _10598_/B _10515_/B vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__a21boi_1
X_13387_ _13386_/A _13386_/B _13386_/C vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15126_ _15433_/CLK _15126_/D _14168_/Y vssd1 vssd1 vccd1 vccd1 _15126_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12338_ _15741_/Q _12339_/B vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15057_ _15107_/CLK _15057_/D _14095_/Y vssd1 vssd1 vccd1 vccd1 _15057_/Q sky130_fd_sc_hd__dfrtp_1
X_12269_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__a21o_1
X_14008_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14008_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater791_A repeater792/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14587__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08500_ _12688_/A vssd1 vssd1 vccd1 vccd1 _08500_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09480_ _09480_/A _09480_/B _09529_/A vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__and3_1
XFILLER_97_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ _08639_/A _08639_/B vssd1 vssd1 vccd1 vccd1 _08666_/A sky130_fd_sc_hd__xnor2_1
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ _15047_/Q vssd1 vssd1 vccd1 vccd1 _13357_/B sky130_fd_sc_hd__buf_6
XFILLER_108_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08293_ _11678_/A vssd1 vssd1 vccd1 vccd1 _08293_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07929__A _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__S _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09816_ _09816_/A _09816_/B _09816_/C vssd1 vssd1 vccd1 vccd1 _09818_/A sky130_fd_sc_hd__and3_1
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09747_ _09747_/A vssd1 vssd1 vccd1 vccd1 _15721_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14497__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11914__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09678_ _15575_/Q vssd1 vssd1 vccd1 vccd1 _09678_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08495__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07695__A1 _07695_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A _08629_/B vssd1 vssd1 vccd1 vccd1 _08629_/X sky130_fd_sc_hd__or2_1
XFILLER_188_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__B_N _15268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11687_/A _11687_/B vssd1 vssd1 vccd1 vccd1 _11642_/C sky130_fd_sc_hd__xnor2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07447__A1 _07447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ _08269_/A _08269_/B _11495_/B _11464_/X vssd1 vssd1 vccd1 vccd1 _11866_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_126_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12745__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13310_/A _13369_/A vssd1 vssd1 vccd1 vccd1 _13312_/B sky130_fd_sc_hd__and2_1
XFILLER_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10522_ _15289_/Q _15256_/Q vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__and2b_1
XFILLER_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _14299_/A vssd1 vssd1 vccd1 vccd1 _14290_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ _10453_/A _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__and3_1
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13241_ _13240_/A _13240_/B _13240_/C vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172_ _13173_/B _13173_/C _13173_/A vssd1 vssd1 vccd1 vccd1 _13247_/B sky130_fd_sc_hd__a21o_2
XANTENNA_input66_A x_i_3[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10383_/A _10383_/C _10383_/B vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__a21oi_1
X_12123_ _12181_/B _12123_/B vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__nand2_2
XFILLER_2_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12054_ _12054_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11005_ _11005_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _15015_/D sky130_fd_sc_hd__nor2_1
XFILLER_133_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15813_ _15813_/A vssd1 vssd1 vccd1 vccd1 _15813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15744_ _15749_/CLK _15744_/D _14821_/Y vssd1 vssd1 vccd1 vccd1 _15744_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14200__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _12956_/A vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__inv_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12639__B _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ _11907_/A vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__inv_2
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15675_ _15707_/CLK _15675_/D _14749_/Y vssd1 vssd1 vccd1 vccd1 _15675_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12887_ _13366_/A _13273_/A vssd1 vssd1 vccd1 vccd1 _12888_/C sky130_fd_sc_hd__xor2_1
XFILLER_209_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _11912_/A _11838_/B vssd1 vssd1 vccd1 vccd1 _11839_/C sky130_fd_sc_hd__and2_1
XFILLER_187_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14557_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14557_/Y sky130_fd_sc_hd__inv_2
X_11769_ _11798_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__xnor2_1
XFILLER_144_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15438_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _13432_/A _13456_/Y _13522_/A vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__mux2_4
XFILLER_173_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14488_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13439_ _13461_/B _13439_/B vssd1 vssd1 vccd1 vccd1 _13441_/C sky130_fd_sc_hd__nand2_1
XFILLER_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater804_A _15586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14870__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08938__A1 _15461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15109_ _15110_/CLK _15109_/D _14150_/Y vssd1 vssd1 vccd1 vccd1 _15109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__A1 _07610_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _15350_/Q _15366_/Q vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__and2b_1
XFILLER_103_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ _09971_/A _07931_/B vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__and2_1
XFILLER_87_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07862_ _15336_/Q input204/X _07900_/S vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09601_ _15425_/Q _15441_/Q vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__or2b_1
XFILLER_113_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07793_ _15370_/Q _07793_/A1 _07803_/S vssd1 vssd1 vccd1 vccd1 _07794_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _15265_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__14110__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07677__A1 _07677_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _15520_/Q _15536_/Q vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__or2b_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ _15049_/Q vssd1 vssd1 vccd1 vccd1 _13422_/A sky130_fd_sc_hd__buf_4
XFILLER_52_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09394_ _09393_/Y _15393_/Q _09392_/B vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__a21o_1
X_08345_ _08324_/A _08324_/B _08344_/X vssd1 vssd1 vccd1 vccd1 _08345_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_196_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08276_ _08325_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_177_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15298__D _15298_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14780__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11909__A _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput460 _15600_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[6] sky130_fd_sc_hd__buf_2
Xoutput471 _11300_/Y vssd1 vssd1 vccd1 vccd1 y_r_4[16] sky130_fd_sc_hd__buf_2
Xoutput482 output482/A vssd1 vssd1 vccd1 vccd1 y_r_5[10] sky130_fd_sc_hd__buf_2
XANTENNA__11628__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput493 output493/A vssd1 vssd1 vccd1 vccd1 y_r_5[5] sky130_fd_sc_hd__buf_2
XFILLER_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15670_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15761__D _15761_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__B _15446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _12810_/A _12810_/B vssd1 vssd1 vccd1 vccd1 _12836_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input120_A x_i_7[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__A0 _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13790_ _13790_/A _13790_/B vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14020__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input218_A x_r_5[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__xor2_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15460_ _15460_/CLK _15460_/D _14522_/Y vssd1 vssd1 vccd1 vccd1 _15460_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _13491_/S _12672_/B vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__nand2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14411_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14411_/Y sky130_fd_sc_hd__inv_2
X_11623_ _11906_/A _12008_/A _11623_/C vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__and3_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15391_/CLK _15391_/D _14449_/Y vssd1 vssd1 vccd1 vccd1 _15391_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_22_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15119_/CLK sky130_fd_sc_hd__clkbuf_16
X_14342_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14342_/Y sky130_fd_sc_hd__inv_2
X_11554_ _11928_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _11623_/C sky130_fd_sc_hd__xor2_2
XFILLER_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _10594_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07840__A1 _07840_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14273_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14273_/Y sky130_fd_sc_hd__inv_2
X_11485_ _08172_/A _08172_/B _11484_/Y vssd1 vssd1 vccd1 vccd1 _11564_/B sky130_fd_sc_hd__a21oi_1
XFILLER_156_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14690__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13224_ _13491_/S _13431_/B _14920_/Q vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__and3_1
XFILLER_170_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _15119_/Q _10296_/Y _10437_/C vssd1 vssd1 vccd1 vccd1 _15809_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11819__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13155_ _13227_/B _12854_/C _13381_/B vssd1 vssd1 vccd1 vccd1 _13156_/B sky130_fd_sc_hd__mux2_1
X_10367_ _10367_/A _10367_/B vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12428_/A _12223_/A _12104_/Y _12105_/Y vssd1 vssd1 vccd1 vccd1 _12152_/A
+ sky130_fd_sc_hd__o31ai_2
XFILLER_111_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07508__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10298_ _15121_/Q _15154_/Q vssd1 vssd1 vccd1 vccd1 _10298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13086_/A _13086_/B vssd1 vssd1 vccd1 vccd1 _13086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output437_A output437/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15363_/CLK sky130_fd_sc_hd__clkbuf_16
X_12037_ _12238_/A vssd1 vssd1 vccd1 vccd1 _12110_/S sky130_fd_sc_hd__inv_2
XFILLER_211_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11554__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13988_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13988_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07659__A1 _07659_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ _15727_/CLK _15727_/D _14804_/Y vssd1 vssd1 vccd1 vccd1 _15727_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _12992_/A _12992_/B vssd1 vssd1 vccd1 vccd1 _12943_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater754_A _15647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14865__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15658_ _15680_/CLK _15658_/D _14731_/Y vssd1 vssd1 vccd1 vccd1 _15658_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14609_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14609_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater921_A input187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ _15725_/CLK _15589_/D _14658_/Y vssd1 vssd1 vccd1 vccd1 _15589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_clk _15044_/CLK vssd1 vssd1 vccd1 vccd1 _15268_/CLK sky130_fd_sc_hd__clkbuf_16
X_08130_ _11707_/A _11617_/A _08144_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__and3_1
XFILLER_109_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08070_/B sky130_fd_sc_hd__xnor2_2
XFILLER_174_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07926__B _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14105__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07418__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08963_ _08963_/A _08963_/B _08963_/C vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__nor3_1
XANTENNA__08103__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _15493_/Q _15477_/Q vssd1 vssd1 vccd1 vccd1 _15218_/D sky130_fd_sc_hd__xor2_1
XFILLER_69_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13944__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08894_ _08957_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _15210_/D sky130_fd_sc_hd__xor2_1
XFILLER_5_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater930 input173/X vssd1 vssd1 vccd1 vccd1 _07828_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07898__A1 input138/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater941 input160/X vssd1 vssd1 vccd1 vccd1 repeater941/X sky130_fd_sc_hd__buf_2
X_07845_ _07845_/A vssd1 vssd1 vccd1 vccd1 _15345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater952 input144/X vssd1 vssd1 vccd1 vccd1 _07886_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater963 input129/X vssd1 vssd1 vccd1 vccd1 _07396_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08996__A_N _15368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__S _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater974 repeater975/X vssd1 vssd1 vccd1 vccd1 _07390_/A1 sky130_fd_sc_hd__buf_4
Xrepeater985 input104/X vssd1 vssd1 vccd1 vccd1 _07514_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_opt_2_0_clk_A _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _07776_/A vssd1 vssd1 vccd1 vccd1 _15379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09515_ _09441_/Y _09514_/B _09443_/B vssd1 vssd1 vccd1 vccd1 _09517_/B sky130_fd_sc_hd__o21ai_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14775__A _14781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09869__A _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09514_/A _09446_/B vssd1 vssd1 vccd1 vccd1 _15275_/D sky130_fd_sc_hd__xor2_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08773__A _15337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09377_ _09377_/A _09377_/B _09377_/C vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__or3_1
XFILLER_184_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08328_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08328_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08075__A1 _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07822__A1 _07822_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _08257_/A _08257_/B _08265_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _15781_/Q vssd1 vssd1 vccd1 vccd1 _11270_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_690 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10709__A1 _15281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10221_ _15075_/Q _15240_/Q vssd1 vssd1 vccd1 vccd1 _10221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14015__A _14017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input168_A x_r_2[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10152_ _10149_/A _10839_/A _10149_/B _10151_/X vssd1 vssd1 vccd1 vccd1 _10155_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput290 output290/A vssd1 vssd1 vccd1 vccd1 y_i_1[6] sky130_fd_sc_hd__buf_2
X_14960_ _15383_/CLK _14960_/D _13992_/Y vssd1 vssd1 vccd1 vccd1 _14960_/Q sky130_fd_sc_hd__dfrtp_1
X_10083_ _15214_/Q _15115_/Q vssd1 vssd1 vccd1 vccd1 _10087_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13911_ _13911_/A _13911_/B vssd1 vssd1 vccd1 vccd1 _15067_/D sky130_fd_sc_hd__xnor2_1
XFILLER_181_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A x_i_1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _15792_/CLK _14891_/D _13920_/Y vssd1 vssd1 vccd1 vccd1 _14891_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11374__A _15752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ _13842_/A _13842_/B _13842_/C vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__or3_1
XFILLER_78_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11093__B _11093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12634__A1 _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ _13783_/B _13772_/B _13772_/C vssd1 vssd1 vccd1 vccd1 _13774_/B sky130_fd_sc_hd__o21a_1
XFILLER_204_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14685__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _15174_/Q vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15512_ _15571_/CLK _15512_/D _14576_/Y vssd1 vssd1 vccd1 vccd1 _15512_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12724_ _12836_/A _12724_/B vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__and2_1
XANTENNA__07510__A0 _15509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08683__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ _15444_/CLK _15443_/D _14504_/Y vssd1 vssd1 vccd1 vccd1 _15443_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_203_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12655_ _12703_/A _12703_/B _12703_/C vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__and3_1
XFILLER_157_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11606_ _11659_/B _11606_/B vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__xnor2_1
XFILLER_180_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15374_ _15374_/CLK _15374_/D _14430_/Y vssd1 vssd1 vccd1 vccd1 _15374_/Q sky130_fd_sc_hd__dfrtp_1
X_12586_ _12586_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _15680_/D sky130_fd_sc_hd__xnor2_1
XFILLER_157_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09802__A2 _15424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output387_A output387/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14325_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14325_/Y sky130_fd_sc_hd__inv_2
X_11537_ _11537_/A _11537_/B _11537_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__and3_1
XFILLER_11_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12933__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14256_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14256_/Y sky130_fd_sc_hd__inv_2
X_11468_ _11832_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15666__D _15666_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _13100_/A _13100_/B _13098_/A _13206_/Y vssd1 vssd1 vccd1 vccd1 _13208_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ _10417_/X _10421_/C vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__and2b_1
X_14187_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07577__A0 _15476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _10207_/Y _11398_/B _10209_/B vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__o21ai_2
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13138_ _13138_/A _13555_/A _13138_/C vssd1 vssd1 vccd1 vccd1 _13213_/A sky130_fd_sc_hd__or3_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13015_/A _13069_/B vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__and2b_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15563_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12873__A1 _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater969_A input122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _15450_/Q input14/X _07632_/S vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _15484_/Q input48/X _07589_/S vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14595__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09300_ _09293_/Y _09298_/B _09295_/B vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__o21ai_1
XFILLER_181_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07492_ _15518_/Q input34/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__mux2_1
XFILLER_185_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ _15497_/Q _15481_/Q vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__and2b_1
XFILLER_179_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09162_ _15566_/Q _15546_/Q vssd1 vssd1 vccd1 vccd1 _09163_/B sky130_fd_sc_hd__nand2_1
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08113_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13939__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _09086_/Y _09091_/B _09088_/B vssd1 vssd1 vccd1 vccd1 _09094_/B sky130_fd_sc_hd__o21ai_1
XFILLER_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08044_ _08045_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__xor2_1
XFILLER_134_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07937__A _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13353__A2 _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09995_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _14932_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08946_ _08862_/Y _08945_/B _08864_/B vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__o21ai_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _08950_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _15207_/D sky130_fd_sc_hd__xor2_2
XFILLER_185_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08487__B _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A _15027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater760 _15642_/Q vssd1 vssd1 vccd1 vccd1 output522/A sky130_fd_sc_hd__clkbuf_2
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _15353_/Q _07828_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07829_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater771 repeater772/X vssd1 vssd1 vccd1 vccd1 output488/A sky130_fd_sc_hd__buf_4
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater782 _15615_/Q vssd1 vssd1 vccd1 vccd1 output493/A sky130_fd_sc_hd__clkbuf_2
Xrepeater793 _15598_/Q vssd1 vssd1 vccd1 vccd1 output458/A sky130_fd_sc_hd__clkbuf_2
X_07759_ _15387_/Q _07759_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07760_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _15719_/Q _15785_/Q vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__and2_1
XFILLER_53_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12737__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09429_ _09504_/A _09426_/B _09428_/X vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__a21o_1
XFILLER_198_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12440_ _12440_/A _12455_/C _12440_/C vssd1 vssd1 vccd1 vccd1 _12463_/B sky130_fd_sc_hd__or3_1
XFILLER_139_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12371_/A _12372_/B _12371_/C vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__nand3_1
XFILLER_154_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _14993_/Q vssd1 vssd1 vccd1 vccd1 _11322_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15090_ _15107_/CLK _15090_/D _14130_/Y vssd1 vssd1 vccd1 vccd1 _15090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14041_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14041_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11253_ _11253_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11253_/Y sky130_fd_sc_hd__nor2_2
XFILLER_84_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07559__A0 _15485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _15071_/Q _10203_/Y _10199_/B vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__a21o_1
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11184_ _15749_/Q _15027_/Q vssd1 vssd1 vccd1 vccd1 _11186_/A sky130_fd_sc_hd__or2_2
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09042__B_N _15377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _15143_/Q _15308_/Q vssd1 vssd1 vccd1 vccd1 _10135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14943_ _15784_/CLK _14943_/D _13974_/Y vssd1 vssd1 vccd1 vccd1 _14943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10066_ _10066_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__nand2_1
XFILLER_208_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12855__A1 _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14874_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14874_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ _13823_/Y _13822_/B _13824_/Y vssd1 vssd1 vccd1 vccd1 _13826_/B sky130_fd_sc_hd__o21ai_2
XFILLER_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output302_A output302/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11832__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13756_ _13848_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _15703_/D sky130_fd_sc_hd__xor2_1
XFILLER_189_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ _10968_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _15006_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12707_ _12945_/A _12930_/A vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13687_ _13684_/A _13822_/A _13686_/Y vssd1 vssd1 vccd1 vccd1 _13696_/A sky130_fd_sc_hd__a21o_1
X_10899_ _14961_/Q _14895_/Q vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15426_ _15438_/CLK _15426_/D _14486_/Y vssd1 vssd1 vccd1 vccd1 _15426_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_549 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12638_ _13203_/A _12945_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ _15719_/CLK _15357_/D _14412_/Y vssd1 vssd1 vccd1 vccd1 _15357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12569_/A _12569_/B vssd1 vssd1 vccd1 vccd1 _15624_/D sky130_fd_sc_hd__xnor2_1
XFILLER_106_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1074 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11594__A1 _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14308_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14308_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15288_ _15542_/CLK _15288_/D _14339_/Y vssd1 vssd1 vccd1 vccd1 _15288_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14239_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14420_/A sky130_fd_sc_hd__buf_8
XFILLER_113_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _15342_/Q _15326_/Q vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__and2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _15432_/Q _15416_/Q _09779_/X vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_674 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08727_/X _08728_/X _08730_/X vssd1 vssd1 vccd1 vccd1 _08731_/X sky130_fd_sc_hd__a21o_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08662_ _08663_/A _08663_/B _08663_/C vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__o21ai_2
XFILLER_187_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07613_ _07613_/A vssd1 vssd1 vccd1 vccd1 _15459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08593_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__and2_1
XFILLER_53_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07544_ _07544_/A vssd1 vssd1 vccd1 vccd1 _15493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07475_ _15526_/Q input90/X _07485_/S vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _15575_/Q _15555_/Q _09213_/X vssd1 vssd1 vccd1 vccd1 _09215_/B sky130_fd_sc_hd__a21oi_2
XFILLER_179_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _15561_/Q _15541_/Q _09628_/C vssd1 vssd1 vccd1 vccd1 _09147_/A sky130_fd_sc_hd__a21oi_1
XFILLER_120_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07789__A0 _15372_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ _09076_/A _09076_/B vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__nor2_2
XFILLER_120_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08047_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _09885_/Y _09977_/B _09887_/B vssd1 vssd1 vccd1 vccd1 _09979_/B sky130_fd_sc_hd__o21ai_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07606__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08929_ _15476_/Q _15460_/Q vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__or2_1
XFILLER_170_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11940_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater590 _10912_/Y vssd1 vssd1 vccd1 vccd1 output309/A sky130_fd_sc_hd__clkbuf_2
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _15732_/Q _11875_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__xnor2_2
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13610_ _13610_/A _13610_/B vssd1 vssd1 vccd1 vccd1 _15094_/D sky130_fd_sc_hd__xor2_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input200_A x_r_4[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822_ _15305_/Q _15140_/Q vssd1 vssd1 vccd1 vccd1 _10823_/C sky130_fd_sc_hd__or2b_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12065__A2 _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14590_ _14600_/A vssd1 vssd1 vccd1 vccd1 _14590_/Y sky130_fd_sc_hd__inv_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09122__A _15504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__nand2_1
XFILLER_198_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _11273_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _10753_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input96_A x_i_5[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ _13428_/A _13428_/B _13426_/A vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__13014__A1 _12945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _10685_/A _11003_/B vssd1 vssd1 vccd1 vccd1 _15047_/D sky130_fd_sc_hd__xor2_4
XFILLER_51_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15211_ _15363_/CLK _15211_/D _14258_/Y vssd1 vssd1 vccd1 vccd1 _15211_/Q sky130_fd_sc_hd__dfrtp_1
X_12423_ _12423_/A _12594_/A _12423_/C vssd1 vssd1 vccd1 vccd1 _12424_/B sky130_fd_sc_hd__nor3_1
XFILLER_205_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ _15406_/CLK _15142_/D _14185_/Y vssd1 vssd1 vccd1 vccd1 _15142_/Q sky130_fd_sc_hd__dfrtp_1
X_12354_ _08347_/A _08347_/B _08347_/C _12353_/X vssd1 vssd1 vccd1 vccd1 _12355_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_181_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _11305_/A _11305_/B vssd1 vssd1 vccd1 vccd1 _11305_/Y sky130_fd_sc_hd__nor2_2
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15073_ _15367_/CLK _15073_/D _14112_/Y vssd1 vssd1 vccd1 vccd1 _15073_/Q sky130_fd_sc_hd__dfrtp_1
X_12285_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__and2_1
XFILLER_142_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08729__C1 _12662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14024_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14024_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11236_ _11235_/A _11235_/B _11385_/A vssd1 vssd1 vccd1 vccd1 _11237_/B sky130_fd_sc_hd__a21oi_2
XFILLER_20_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11167_ _11167_/A _11359_/A _11167_/C vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__and3_1
XFILLER_96_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14203__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ _10112_/A _10114_/B _10112_/B vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__11546__B _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ _15002_/Q _14936_/Q vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__and2b_1
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output517_A output517/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09016__B _15356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10049_ _10043_/A _10045_/B _10043_/B vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__a21boi_2
X_14926_ _15221_/CLK _14926_/D _13956_/Y vssd1 vssd1 vccd1 vccd1 _14926_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14857_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14857_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater667_A _14737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15044__CLK _15044_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ _13808_/A _14938_/Q vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__or2b_2
XFILLER_95_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14788_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14788_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13739_ _13740_/B _13740_/C _13740_/A vssd1 vssd1 vccd1 vccd1 _13741_/A sky130_fd_sc_hd__a21oi_1
XFILLER_56_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater834_A input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14873__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ _15588_/CLK _15409_/D _14468_/Y vssd1 vssd1 vccd1 vccd1 _15409_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_83_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09901_ _15191_/Q _15224_/Q vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09832_ _09832_/A _09832_/B _09832_/C vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__and3_1
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07934__B _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10641__A _15270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12819__A1 _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _15067_/Q _15100_/Q _09762_/B vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__a21oi_2
XFILLER_101_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13952__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _08631_/X _08633_/A _08713_/Y vssd1 vssd1 vccd1 vccd1 _08714_/X sky130_fd_sc_hd__a21bo_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09694_ _15056_/Q _15089_/Q vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__or2_1
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _12945_/A _12881_/A _08645_/C vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__and3_1
XFILLER_82_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ _08629_/A _08629_/B _08551_/A vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__a21bo_1
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11191__B _15028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _07527_/A vssd1 vssd1 vccd1 vccd1 _15501_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14783__A _14784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07458_ _07458_/A vssd1 vssd1 vccd1 vccd1 _15535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07389_ _07389_/A vssd1 vssd1 vccd1 vccd1 _15573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ _15506_/Q _15490_/Q vssd1 vssd1 vccd1 vccd1 _09265_/A sky130_fd_sc_hd__xnor2_2
XFILLER_135_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ _15380_/Q _15364_/Q vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__nand2_1
XFILLER_194_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _12254_/A vssd1 vssd1 vccd1 vccd1 _12132_/S sky130_fd_sc_hd__inv_2
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11647__A _12378_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ _14987_/Q _11021_/B vssd1 vssd1 vccd1 vccd1 _11021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input150_A x_r_1[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14023__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input248_A x_r_7[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08021__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _15761_/CLK _15760_/D _14838_/Y vssd1 vssd1 vccd1 vccd1 _15760_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12874_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__and2b_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_715 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A x_i_0[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _11846_/A _11846_/B _11922_/X vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__a21oi_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14714_/A vssd1 vssd1 vccd1 vccd1 _14711_/Y sky130_fd_sc_hd__inv_2
X_15691_ _15699_/CLK _15691_/D _14766_/Y vssd1 vssd1 vccd1 vccd1 _15691_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__buf_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _11855_/A _11855_/B _11855_/C vssd1 vssd1 vccd1 vccd1 _11931_/A sky130_fd_sc_hd__a21o_1
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_972 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10805_ _15725_/Q _15791_/Q vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14573_/Y sky130_fd_sc_hd__inv_2
X_11785_ _11787_/B _11787_/C vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__and2_1
XANTENNA__14693__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13524_ _13524_/A _13524_/B vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__xnor2_2
XFILLER_201_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10736_ _10734_/Y _10736_/B vssd1 vssd1 vccd1 vccd1 _11259_/A sky130_fd_sc_hd__and2b_1
XFILLER_201_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14904__CLK _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12925__B _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13455_ _13455_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__nand2_1
XFILLER_201_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10667_ _10665_/Y _10667_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__and2b_1
XFILLER_16_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12406_ _12406_/A _12406_/B _12406_/C vssd1 vssd1 vccd1 vccd1 _12407_/B sky130_fd_sc_hd__and3_1
XFILLER_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13386_ _13386_/A _13386_/B _13386_/C vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__and3_1
XFILLER_63_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10598_ _10598_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _14992_/D sky130_fd_sc_hd__xnor2_1
XFILLER_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output467_A output467/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ _15433_/CLK _15125_/D _14167_/Y vssd1 vssd1 vccd1 vccd1 _15125_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12337_ _12520_/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12339_/B sky130_fd_sc_hd__xnor2_2
XFILLER_103_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15056_ _15712_/CLK _15056_/D _14094_/Y vssd1 vssd1 vccd1 vccd1 _15056_/Q sky130_fd_sc_hd__dfrtp_1
X_12268_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__and3_1
XFILLER_123_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14007_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14007_/Y sky130_fd_sc_hd__inv_2
X_11219_ _11219_/A vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12199_ _12252_/B _12199_/B vssd1 vssd1 vccd1 vccd1 _12201_/C sky130_fd_sc_hd__or2_1
XFILLER_122_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater784_A _15608_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14868__A _14872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput190 x_r_3[5] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _15528_/CLK _14909_/D _13939_/Y vssd1 vssd1 vccd1 vccd1 _14909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ _08663_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08639_/B sky130_fd_sc_hd__and2b_1
XFILLER_184_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _08728_/B _08369_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__or3b_1
XFILLER_189_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ _11832_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08292_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_176_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07929__B _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10636__A _15269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14108__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13012__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13947__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12851__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11467__A _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1002 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input3_A x_i_0[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _15053_/Q _09687_/Y _09816_/C vssd1 vssd1 vccd1 vccd1 _15743_/D sky130_fd_sc_hd__o21a_1
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14778__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__A1 _07392_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09746_ _09744_/X _09752_/A vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__and2b_1
XFILLER_189_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11206__B_N _15030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A _09677_/B vssd1 vssd1 vccd1 vccd1 _15314_/D sky130_fd_sc_hd__nor2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ _08716_/A _08718_/B _08627_/X vssd1 vssd1 vccd1 vccd1 _08633_/B sky130_fd_sc_hd__o21ai_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _13145_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _08560_/B sky130_fd_sc_hd__or2_1
XFILLER_196_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11865_/C sky130_fd_sc_hd__nor2_1
XFILLER_168_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1085 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12745__B _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15759__D _15759_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_805 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _10519_/Y _10521_/B vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__nand2b_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input198_A x_r_4[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14018__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ _13240_/A _13240_/B _13240_/C vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__and3_1
XFILLER_202_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10452_ _15157_/Q _15124_/Q vssd1 vssd1 vccd1 vccd1 _10453_/C sky130_fd_sc_hd__or2b_1
XFILLER_182_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _13247_/A _13171_/B vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__nand2_1
X_10383_ _10383_/A _10383_/B _10383_/C vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__and3_1
X_12122_ _12122_/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__or2_1
XANTENNA__13576__B _13576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A x_i_3[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12053_ _12053_/A _12053_/B _12053_/C vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__and3_1
XFILLER_46_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11003_/A _11003_/C _11003_/B vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__a21oi_1
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14688__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15812_ _15812_/A vssd1 vssd1 vccd1 vccd1 _15812_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13456__A1 _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15743_ _15777_/CLK _15743_/D _14820_/Y vssd1 vssd1 vccd1 vccd1 _15743_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _13116_/B _12955_/B vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11906_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__nand2_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12886_/A vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__inv_2
X_15674_ _15707_/CLK _15674_/D _14748_/Y vssd1 vssd1 vccd1 vccd1 _15674_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _12312_/S _12204_/A vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__or2_1
X_14625_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14625_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14556_/Y sky130_fd_sc_hd__inv_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11799_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10719_ _15710_/Q _15776_/Q vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__or2b_1
X_13507_ _13490_/A _13490_/B _13492_/B vssd1 vssd1 vccd1 vccd1 _13522_/A sky130_fd_sc_hd__o21ai_1
XFILLER_13_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater532_A _12221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14487_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ _11740_/A _11478_/B _11906_/A vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__mux2_1
XFILLER_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13438_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13439_/B sky130_fd_sc_hd__or2_1
XFILLER_173_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08938__A2 _15445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ _13369_/A _13369_/B _13369_/C vssd1 vssd1 vccd1 vccd1 _13370_/B sky130_fd_sc_hd__and3_1
XFILLER_6_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _15750_/CLK _15108_/D _14149_/Y vssd1 vssd1 vccd1 vccd1 _15108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07930_ _15185_/Q _15218_/Q vssd1 vssd1 vccd1 vccd1 _07931_/B sky130_fd_sc_hd__or2_1
X_15039_ _15525_/CLK _15039_/D _14076_/Y vssd1 vssd1 vccd1 vccd1 _15039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10191__A _15218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07861_ _07861_/A vssd1 vssd1 vccd1 vccd1 _15337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15382__CLK _15666_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14598__A _14600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _15179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07792_ _07792_/A vssd1 vssd1 vccd1 vccd1 _15371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07704__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ _09529_/A _09529_/B _09530_/X vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09462_ _09462_/A vssd1 vssd1 vccd1 vccd1 _15277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08413_ _13366_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09393_ _15409_/Q vssd1 vssd1 vccd1 vccd1 _09393_/Y sky130_fd_sc_hd__inv_2
X_08344_ _08325_/X _08277_/Y _08343_/X vssd1 vssd1 vccd1 vccd1 _08344_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08275_ _08322_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13677__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1007 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11909__B _12247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput450 output450/A vssd1 vssd1 vccd1 vccd1 y_r_3[12] sky130_fd_sc_hd__buf_2
Xoutput461 output461/A vssd1 vssd1 vccd1 vccd1 y_r_3[7] sky130_fd_sc_hd__buf_2
XFILLER_191_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput472 output472/A vssd1 vssd1 vccd1 vccd1 y_r_4[1] sky130_fd_sc_hd__buf_2
Xoutput483 _15621_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[11] sky130_fd_sc_hd__buf_2
XFILLER_121_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput494 output494/A vssd1 vssd1 vccd1 vccd1 y_r_5[6] sky130_fd_sc_hd__buf_2
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14301__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09729_ _15063_/Q _15096_/Q vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__or2b_1
XFILLER_170_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _12871_/A _08520_/C _12739_/Y vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_input113_A x_i_6[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A _12735_/C vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__xnor2_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14410_ _14419_/A vssd1 vssd1 vccd1 vccd1 _14410_/Y sky130_fd_sc_hd__inv_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11622_/A _11707_/A _11687_/A vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__and3_1
XFILLER_169_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15390_ _15391_/CLK _15390_/D _14448_/Y vssd1 vssd1 vccd1 vccd1 _15390_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _14359_/A vssd1 vssd1 vccd1 vccd1 _14341_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11553_ _11906_/A _12008_/A vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__nand2_1
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ _10594_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _15023_/D sky130_fd_sc_hd__xor2_1
X_14272_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14272_/Y sky130_fd_sc_hd__inv_2
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11484_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _13431_/B _13223_/B vssd1 vssd1 vccd1 vccd1 _13320_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10435_ _10104_/Y _15152_/Q _10296_/B vssd1 vssd1 vccd1 vccd1 _10437_/C sky130_fd_sc_hd__a21o_1
XFILLER_124_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13913__A2 _15331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ _13390_/A vssd1 vssd1 vccd1 vccd1 _13227_/B sky130_fd_sc_hd__inv_2
XFILLER_83_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10366_ _15166_/Q _15133_/Q vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__and2b_1
XFILLER_88_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12105_ _12451_/B _12105_/B vssd1 vssd1 vccd1 vccd1 _12105_/Y sky130_fd_sc_hd__nand2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13085_ _13175_/A _13175_/B vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__xnor2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10297_ _15120_/Q _15153_/Q _10296_/Y _10104_/Y vssd1 vssd1 vccd1 vccd1 _10301_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12036_ _12038_/A _12122_/A _12231_/A _11956_/X _12238_/A vssd1 vssd1 vccd1 vccd1
+ _12040_/A sky130_fd_sc_hd__o2111a_1
XANTENNA__13141__A3 _13713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output332_A _11346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14211__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__B _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13987_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13987_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15726_ _15727_/CLK _15726_/D _14803_/Y vssd1 vssd1 vccd1 vccd1 _15726_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _13012_/A _12892_/B _12896_/B _12937_/Y vssd1 vssd1 vccd1 vccd1 _12992_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15657_ _15784_/CLK _15657_/D _14730_/Y vssd1 vssd1 vccd1 vccd1 _15657_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater747_A repeater748/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12869_ _12798_/A _12798_/B _12868_/X vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__12666__A _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__B _15449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14608_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15588_ _15588_/CLK _15588_/D _14657_/Y vssd1 vssd1 vccd1 vccd1 _15588_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14539_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14539_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater914_A input199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14881__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08962_ _15471_/Q _15455_/Q vssd1 vssd1 vccd1 vccd1 _08963_/C sky130_fd_sc_hd__and2_1
XFILLER_9_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07913_ _07913_/A vssd1 vssd1 vccd1 vccd1 _15086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08893_ _08955_/A _08887_/B _08892_/X vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__a21o_1
XFILLER_124_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater920 input188/X vssd1 vssd1 vccd1 vccd1 _07700_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater931 input172/X vssd1 vssd1 vccd1 vccd1 _07830_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07942__B _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07844_ _15345_/Q _07844_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14121__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater942 input159/X vssd1 vssd1 vccd1 vccd1 _07759_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater953 input143/X vssd1 vssd1 vccd1 vccd1 _07888_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_151_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater964 input128/X vssd1 vssd1 vccd1 vccd1 _07398_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater975 input117/X vssd1 vssd1 vccd1 vccd1 repeater975/X sky130_fd_sc_hd__buf_2
XFILLER_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater986 input103/X vssd1 vssd1 vccd1 vccd1 _07516_/A1 sky130_fd_sc_hd__clkbuf_2
X_07775_ _15379_/Q input232/X _07803_/S vssd1 vssd1 vccd1 vccd1 _07776_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13960__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _15259_/D sky130_fd_sc_hd__xor2_1
XFILLER_140_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _09511_/A _09440_/B _09444_/X vssd1 vssd1 vccd1 vccd1 _09446_/B sky130_fd_sc_hd__a21o_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12576__A _14939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08773__B _15321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09376_ _15405_/Q _15389_/Q vssd1 vssd1 vccd1 vccd1 _09377_/C sky130_fd_sc_hd__and2b_1
XFILLER_36_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08327_/X sky130_fd_sc_hd__and2_1
XFILLER_184_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08075__A2 _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14791__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _08281_/A _08281_/B vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14941__D _14941_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _08189_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13200__A _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _11400_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__nand2_1
XFILLER_180_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10151_ _15145_/Q _15310_/Q vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__and2_1
XFILLER_161_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput280 output280/A vssd1 vssd1 vccd1 vccd1 y_i_1[12] sky130_fd_sc_hd__buf_2
XFILLER_0_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput291 _15650_/Q vssd1 vssd1 vccd1 vccd1 y_i_1[7] sky130_fd_sc_hd__buf_2
XFILLER_88_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ _10082_/A vssd1 vssd1 vccd1 vccd1 _14983_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input230_A x_r_6[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13910_ _13908_/A _13908_/B _13909_/X vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__a21o_1
X_14890_ _15809_/CLK _14890_/D _13919_/Y vssd1 vssd1 vccd1 vccd1 _14890_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14031__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11374__B _15030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _13841_/A _13841_/B _14979_/Q vssd1 vssd1 vccd1 vccd1 _13842_/C sky130_fd_sc_hd__nor3b_1
XFILLER_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13870__A _14985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ _13783_/B _13772_/B _13772_/C vssd1 vssd1 vccd1 vccd1 _13774_/A sky130_fd_sc_hd__nor3_1
XFILLER_210_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10984_ _10984_/A _10984_/B vssd1 vssd1 vccd1 vccd1 _15010_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15511_ _15511_/CLK _15511_/D _14575_/Y vssd1 vssd1 vccd1 vccd1 _15511_/Q sky130_fd_sc_hd__dfrtp_4
X_12723_ _12723_/A _12726_/A _12723_/C vssd1 vssd1 vccd1 vccd1 _12724_/B sky130_fd_sc_hd__or3_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07510__A1 _07510_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__S _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15442_ _15732_/CLK _15442_/D _14503_/Y vssd1 vssd1 vccd1 vccd1 _15442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12703_/C sky130_fd_sc_hd__xnor2_1
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11605_ _11526_/A _11526_/B _11604_/Y vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _12585_/A _12585_/B vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__nand2_1
X_15373_ _15617_/CLK _15373_/D _14429_/Y vssd1 vssd1 vccd1 vccd1 _15373_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ _11537_/A _11537_/B _11537_/C vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__a21oi_1
X_14324_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14324_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output282_A output282/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14255_/Y sky130_fd_sc_hd__inv_2
X_11467_ _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14206__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13110__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ _13206_/A vssd1 vssd1 vccd1 vccd1 _13206_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ _10417_/B _10417_/C _10417_/A vssd1 vssd1 vccd1 vccd1 _10421_/C sky130_fd_sc_hd__a21o_1
X_14186_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14186_/Y sky130_fd_sc_hd__inv_2
X_11398_ _11398_/A _11398_/B vssd1 vssd1 vccd1 vccd1 _15730_/D sky130_fd_sc_hd__xnor2_1
XFILLER_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07577__A1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13555_/A _13137_/B vssd1 vssd1 vccd1 vccd1 _15633_/D sky130_fd_sc_hd__xor2_1
X_10349_ _15131_/Q _15164_/Q vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__and2b_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A _13552_/A vssd1 vssd1 vccd1 vccd1 _15632_/D sky130_fd_sc_hd__xor2_1
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15682__D _15682_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater697_A _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08858__B _15448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _12223_/A _12223_/B vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_420 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14876__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater864_A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07560_ _07560_/A vssd1 vssd1 vccd1 vccd1 _15485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15709_ _15777_/CLK _15709_/D _14785_/Y vssd1 vssd1 vccd1 vccd1 _15709_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07491_ _07491_/A vssd1 vssd1 vccd1 vccd1 _15519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ _09230_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _15238_/D sky130_fd_sc_hd__xor2_2
XFILLER_94_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_827 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09161_ _15566_/Q _15546_/Q vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08112_ _08112_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__xnor2_1
XFILLER_175_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _15499_/Q _15483_/Q vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__xnor2_2
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__xnor2_1
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14116__A _14118_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1135 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13955__A _13957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_992 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09994_ _09993_/B _09993_/C _09993_/A vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__o21a_1
XFILLER_89_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _15189_/D sky130_fd_sc_hd__xor2_1
XFILLER_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15592__D _15592_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08876_ _08947_/A _08871_/B _08875_/X vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__a21o_1
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater750 _15652_/Q vssd1 vssd1 vccd1 vccd1 output293/A sky130_fd_sc_hd__clkbuf_2
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _07827_/A vssd1 vssd1 vccd1 vccd1 _15354_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater761 _15641_/Q vssd1 vssd1 vccd1 vccd1 output521/A sky130_fd_sc_hd__clkbuf_2
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater772 _15626_/Q vssd1 vssd1 vccd1 vccd1 repeater772/X sky130_fd_sc_hd__buf_2
XFILLER_178_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07740__A1 _07740_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater783 _15609_/Q vssd1 vssd1 vccd1 vccd1 output453/A sky130_fd_sc_hd__buf_4
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater794 _15595_/Q vssd1 vssd1 vccd1 vccd1 output455/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07758_ _07758_/A vssd1 vssd1 vccd1 vccd1 _15388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08296__A2 _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07689_ _15421_/Q _07689_/A1 _07695_/S vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12737__C _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09428_ _15529_/Q _15513_/Q vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__and2b_1
XFILLER_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ _09359_/A _09359_/B vssd1 vssd1 vccd1 vccd1 _15138_/D sky130_fd_sc_hd__xor2_1
XFILLER_8_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08008__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12370_ _12371_/A _12371_/C _12372_/B _12372_/A vssd1 vssd1 vccd1 vccd1 _12373_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input180_A x_r_3[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14026__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ _14058_/A vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__inv_2
X_11252_ _11251_/A _11251_/C _11251_/B vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__a21oi_1
XFILLER_153_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11369__B _11369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07559__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _15236_/Q vssd1 vssd1 vccd1 vccd1 _10203_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11183_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input41_A x_i_2[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _10828_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _15799_/D sky130_fd_sc_hd__xnor2_1
XFILLER_171_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_916 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14942_ _15732_/CLK _14942_/D _13973_/Y vssd1 vssd1 vccd1 vccd1 _14942_/Q sky130_fd_sc_hd__dfrtp_1
X_10065_ _10066_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _14981_/D sky130_fd_sc_hd__xor2_2
XANTENNA__12855__A2 _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14873_ _14881_/A vssd1 vssd1 vccd1 vccd1 _14873_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14696__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _14975_/Q _13824_/B vssd1 vssd1 vccd1 vccd1 _13824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10967_ _10966_/A _10966_/C _10966_/B vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__a21oi_1
X_13755_ _13743_/A _13842_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__o21a_1
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _13203_/A _12813_/C vssd1 vssd1 vccd1 vccd1 _12930_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10898_ _14961_/Q _14895_/Q vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__or2_1
X_13686_ _13686_/A _13824_/B vssd1 vssd1 vccd1 vccd1 _13686_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_output497_A _15619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15425_ _15438_/CLK _15425_/D _14485_/Y vssd1 vssd1 vccd1 vccd1 _15425_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _13352_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ _12567_/Y _12566_/B _12298_/A vssd1 vssd1 vccd1 vccd1 _12569_/B sky130_fd_sc_hd__a21oi_1
X_15356_ _15758_/CLK _15356_/D _14411_/Y vssd1 vssd1 vccd1 vccd1 _15356_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15677__D _15677_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ _12231_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14307_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12499_ _12610_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _15656_/D sky130_fd_sc_hd__xnor2_1
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15287_ _15592_/CLK _15287_/D _14338_/Y vssd1 vssd1 vccd1 vccd1 _15287_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14238_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14238_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14169_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14169_/Y sky130_fd_sc_hd__inv_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _12654_/A _12688_/A _08726_/Y _08729_/X vssd1 vssd1 vccd1 vccd1 _08730_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08661_ _08661_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _08663_/C sky130_fd_sc_hd__xnor2_1
XFILLER_38_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07722__A1 _07722_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07612_ _15459_/Q input8/X _07632_/S vssd1 vssd1 vccd1 vccd1 _07613_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08592_ _08592_/A _08594_/A vssd1 vssd1 vccd1 vccd1 _08633_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07543_ _15493_/Q _07543_/A1 _07591_/S vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__mux2_1
XFILLER_207_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07474_ _07474_/A vssd1 vssd1 vccd1 vccd1 _15527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ _15575_/Q _15555_/Q _09208_/A vssd1 vssd1 vccd1 vccd1 _09213_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12854__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09144_ _09631_/A _09144_/B vssd1 vssd1 vccd1 vccd1 _09628_/C sky130_fd_sc_hd__nand2_1
XFILLER_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_775 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07789__A1 _07789_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _15495_/Q _15479_/Q vssd1 vssd1 vccd1 vccd1 _09076_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08026_ _08026_/A _08025_/X vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__or2b_1
XFILLER_151_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08779__A _15338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07410__A0 _15562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09977_ _09977_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _14925_/D sky130_fd_sc_hd__xnor2_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _15476_/Q _15460_/Q vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _15463_/Q vssd1 vssd1 vccd1 vccd1 _08859_/Y sky130_fd_sc_hd__inv_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater580 repeater581/X vssd1 vssd1 vccd1 vccd1 output343/A sky130_fd_sc_hd__buf_4
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11870_/A _12406_/A vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__xor2_2
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater591 _11324_/X vssd1 vssd1 vccd1 vccd1 output342/A sky130_fd_sc_hd__clkbuf_2
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07622__S _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10823_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10487__B_N _15252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10549__A _15294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _10744_/Y _10748_/B _10746_/B vssd1 vssd1 vccd1 vccd1 _10753_/B sky130_fd_sc_hd__o21ai_2
X_13540_ _13538_/Y _13536_/A _13536_/B _13539_/Y vssd1 vssd1 vccd1 vccd1 _13541_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09122__B _15488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08019__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13471_ _13471_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__nor2_2
XFILLER_201_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10683_ _15278_/Q _15179_/Q vssd1 vssd1 vccd1 vccd1 _11003_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09218__A1 _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12422_ _12423_/A _12423_/C _12594_/A vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__o21a_1
X_15210_ _15363_/CLK _15210_/D _14257_/Y vssd1 vssd1 vccd1 vccd1 _15210_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input89_A x_i_5[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ _11499_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__and2b_1
XFILLER_154_723 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15141_ _15406_/CLK _15141_/D _14184_/Y vssd1 vssd1 vccd1 vccd1 _15141_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11304_ _11303_/A _11303_/C _11303_/B vssd1 vssd1 vccd1 vccd1 _11305_/B sky130_fd_sc_hd__a21oi_1
X_15072_ _15712_/CLK _15072_/D _14111_/Y vssd1 vssd1 vccd1 vccd1 _15072_/Q sky130_fd_sc_hd__dfrtp_1
X_12284_ _12284_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14023_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14023_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08729__B1 _12627_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11235_ _11235_/A _11235_/B _11385_/A vssd1 vssd1 vccd1 vccd1 _11237_/A sky130_fd_sc_hd__and3_1
XFILLER_153_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07593__A _07805_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11166_ _15023_/Q _15745_/Q vssd1 vssd1 vccd1 vccd1 _11167_/C sky130_fd_sc_hd__or2b_1
XFILLER_121_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10117_ _10115_/Y _10117_/B vssd1 vssd1 vccd1 vccd1 _10817_/A sky130_fd_sc_hd__nand2b_1
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ _14936_/Q _15002_/Q vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__and2b_1
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _15220_/CLK _14925_/D _13955_/Y vssd1 vssd1 vccd1 vccd1 _14925_/Q sky130_fd_sc_hd__dfrtp_1
X_10048_ _10046_/Y _10048_/B vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__and2b_1
XANTENNA_output412_A output412/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07704__A1 _07704_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_784 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11843__A _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14856_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07532__S _07532_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13807_ _13807_/A _13873_/A vssd1 vssd1 vccd1 vccd1 _15708_/D sky130_fd_sc_hd__xnor2_1
XFILLER_63_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater562_A _11285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14787_ _14787_/A vssd1 vssd1 vccd1 vccd1 _14787_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11999_ _11999_/A _11999_/B vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__and2_1
XFILLER_1_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_664 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13738_ _13744_/A _13744_/B vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__xnor2_1
XFILLER_91_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12674__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ _13669_/A _13669_/B vssd1 vssd1 vccd1 vccd1 _13669_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_repeater827_A input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_807 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15408_ _15588_/CLK _15408_/D _14467_/Y vssd1 vssd1 vccd1 vccd1 _15408_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _15374_/CLK _15339_/D _14393_/Y vssd1 vssd1 vccd1 vccd1 _15339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07640__A0 _15445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09900_ _15191_/Q _15224_/Q vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09831_ _15091_/Q _15058_/Q vssd1 vssd1 vccd1 vccd1 _09832_/C sky130_fd_sc_hd__or2b_1
XFILLER_28_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09762_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _15723_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08713_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08713_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09693_ _09693_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _15711_/D sky130_fd_sc_hd__xnor2_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08644_ _12810_/A _08644_/B vssd1 vssd1 vccd1 vccd1 _08649_/A sky130_fd_sc_hd__nor2_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08575_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08631_/A sky130_fd_sc_hd__or2_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07526_ _15501_/Q _07526_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__mux2_1
XFILLER_211_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_887 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ _15535_/Q _07457_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11007__A1 _15278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13399__B _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ _15573_/Q _07388_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07389_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _09125_/A _09258_/B _09126_/X vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__a21oi_1
XFILLER_210_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _15116_/D sky130_fd_sc_hd__nor2_1
XFILLER_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08009_ _11797_/A _11658_/A _08009_/C vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__and3_1
XANTENNA__11928__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14304__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11020_/A _11021_/B vssd1 vssd1 vccd1 vccd1 _11020_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input143_A x_r_0[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _13054_/A _13054_/B vssd1 vssd1 vccd1 vccd1 _13052_/B sky130_fd_sc_hd__xor2_4
XANTENNA__15780__D _15780_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11663__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14710_/Y sky130_fd_sc_hd__inv_2
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11845_/B _11922_/B vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__and2b_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_727 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15690_ _15690_/CLK _15690_/D _14765_/Y vssd1 vssd1 vccd1 vccd1 _15690_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14842_/A vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__buf_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11855_/C sky130_fd_sc_hd__nand2_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _10802_/A _11298_/A _10803_/Y vssd1 vssd1 vccd1 vccd1 _10806_/A sky130_fd_sc_hd__o21ai_1
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11784_ _11783_/A _11783_/B _12391_/B vssd1 vssd1 vccd1 vccd1 _11787_/C sky130_fd_sc_hd__o21bai_1
X_14572_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14572_/Y sky130_fd_sc_hd__inv_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13431_/B _13522_/Y _14920_/Q vssd1 vssd1 vccd1 vccd1 _13524_/B sky130_fd_sc_hd__o21a_2
X_10735_ _15713_/Q _15779_/Q vssd1 vssd1 vccd1 vccd1 _10736_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07870__A0 _15332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10666_ _15275_/Q _15176_/Q vssd1 vssd1 vccd1 vccd1 _10667_/B sky130_fd_sc_hd__nand2_1
X_13454_ _13448_/A _13769_/B _13453_/X vssd1 vssd1 vccd1 vccd1 _13475_/A sky130_fd_sc_hd__a21bo_1
XFILLER_127_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ _12406_/B _12406_/C _12406_/A vssd1 vssd1 vccd1 vccd1 _12455_/D sky130_fd_sc_hd__a21oi_2
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13385_ _13385_/A _13385_/B vssd1 vssd1 vccd1 vccd1 _13386_/C sky130_fd_sc_hd__or2_1
XFILLER_16_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10597_ _10506_/Y _10596_/B _10508_/B vssd1 vssd1 vccd1 vccd1 _10598_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15020__D _15020_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15433_/CLK _15124_/D _14166_/Y vssd1 vssd1 vccd1 vccd1 _15124_/Q sky130_fd_sc_hd__dfrtp_1
X_12336_ _12334_/Y _12317_/B _12335_/Y vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__a21oi_2
XFILLER_154_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12267_ _12563_/A vssd1 vssd1 vccd1 vccd1 _12268_/C sky130_fd_sc_hd__inv_2
X_15055_ _15352_/CLK _15055_/D _14093_/Y vssd1 vssd1 vccd1 vccd1 _15055_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14214__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14006_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14006_/Y sky130_fd_sc_hd__inv_2
X_11218_ _11216_/X _11223_/B vssd1 vssd1 vccd1 vccd1 _11218_/X sky130_fd_sc_hd__and2b_1
XFILLER_96_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ _12197_/B _12198_/B vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__and2b_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11149_ _15709_/Q _11147_/Y _11153_/B vssd1 vssd1 vccd1 vccd1 _11149_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput180 x_r_3[10] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_hd__clkbuf_2
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput191 x_r_3[6] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14908_ _15399_/CLK _14908_/D _13937_/Y vssd1 vssd1 vccd1 vccd1 _14908_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09043__A _15377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14839_ _14841_/A vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14884__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _12881_/A _12654_/A vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__xor2_2
XFILLER_108_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14124__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07437__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09814_ _09688_/Y _15086_/Q _09687_/B vssd1 vssd1 vccd1 vccd1 _09816_/C sky130_fd_sc_hd__a21o_1
XFILLER_115_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13963__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07961__A _15152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09745_ _09744_/A _09744_/B _09857_/A vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09675_/A _09675_/C _09675_/B vssd1 vssd1 vccd1 vccd1 _09677_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_979 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08716_/A _08718_/B _08601_/X _08626_/X vssd1 vssd1 vccd1 vccd1 _08627_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14794__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08558_ _08558_/A _08567_/A vssd1 vssd1 vccd1 vccd1 _08629_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07900__S _07900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14944__D _14944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ _07509_/A vssd1 vssd1 vccd1 vccd1 _15510_/D sky130_fd_sc_hd__clkbuf_1
X_08489_ _08728_/A _12662_/A _08488_/X _08552_/A vssd1 vssd1 vccd1 vccd1 _08548_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13203__A _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ _15257_/Q _15290_/Q vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__nand2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_817 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10451_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10453_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07604__A0 _15463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _13170_/A _13170_/B _13168_/Y vssd1 vssd1 vccd1 vccd1 _13171_/B sky130_fd_sc_hd__or3b_1
X_10382_ _07939_/A _10380_/Y _10383_/C vssd1 vssd1 vccd1 vccd1 _14939_/D sky130_fd_sc_hd__o21a_1
X_12121_ _12122_/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12181_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11658__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14034__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _12053_/A _12053_/B _12053_/C vssd1 vssd1 vccd1 vccd1 _12054_/A sky130_fd_sc_hd__a21oi_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11003_ _11003_/A _11003_/B _11003_/C vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__and3_1
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15811_ _15811_/A vssd1 vssd1 vccd1 vccd1 _15811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15742_ _15791_/CLK _15742_/D _14819_/Y vssd1 vssd1 vccd1 vccd1 _15742_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_82_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _13390_/A _13319_/A _12953_/C vssd1 vssd1 vccd1 vccd1 _12955_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08332__A1 _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11905_ _11905_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__xor2_4
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15673_ _15708_/CLK _15673_/D _14747_/Y vssd1 vssd1 vccd1 vccd1 _15673_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12824_/S _12921_/A _12881_/A _12825_/A _12884_/X vssd1 vssd1 vccd1 vccd1
+ _12886_/A sky130_fd_sc_hd__a41o_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14624_/Y sky130_fd_sc_hd__inv_2
X_11836_ _12312_/S _12204_/A vssd1 vssd1 vccd1 vccd1 _11912_/A sky130_fd_sc_hd__nand2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07810__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_97_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_662 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14555_/Y sky130_fd_sc_hd__inv_2
X_11767_ _11767_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__xnor2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14209__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13506_ _13417_/B _13504_/X _13506_/S vssd1 vssd1 vccd1 vccd1 _13803_/A sky130_fd_sc_hd__mux2_2
XFILLER_187_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ _15776_/Q _15710_/Q vssd1 vssd1 vccd1 vccd1 _11251_/A sky130_fd_sc_hd__or2b_1
XFILLER_201_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14486_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14486_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11698_ _11928_/A vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_20_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__nand2_1
X_10649_ _10974_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _15040_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__12952__A _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12195__A2 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _13369_/A _13369_/B _13369_/C vssd1 vssd1 vccd1 vccd1 _13370_/A sky130_fd_sc_hd__a21oi_1
XFILLER_138_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15107_ _15107_/CLK _15107_/D _14148_/Y vssd1 vssd1 vccd1 vccd1 _15107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12319_ _12319_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__and2_1
X_13299_ _13422_/A _13366_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13300_/B sky130_fd_sc_hd__and3b_1
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ _15509_/CLK _15038_/D _14075_/Y vssd1 vssd1 vccd1 vccd1 _15038_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater894_A input228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14879__A _14881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ _15337_/Q input205/X _07892_/S vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07791_ _15371_/Q input239/X _07791_/S vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _15538_/Q _15522_/Q vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__and2_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09461_ _09459_/X _09466_/B vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__and2b_1
XFILLER_37_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _08412_/A _08412_/B vssd1 vssd1 vccd1 vccd1 _08429_/B sky130_fd_sc_hd__and2_1
XFILLER_184_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09392_/A _09392_/B vssd1 vssd1 vccd1 vccd1 _15147_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10548__B_N _15294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _08325_/X _08277_/Y _08326_/X _08341_/X _08342_/X vssd1 vssd1 vccd1 vccd1
+ _08343_/X sky130_fd_sc_hd__o221a_1
XFILLER_178_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14119__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08274_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__xor2_1
XFILLER_177_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08117__A _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13958__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11478__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput440 output440/A vssd1 vssd1 vccd1 vccd1 y_r_2[3] sky130_fd_sc_hd__buf_2
Xoutput451 output451/A vssd1 vssd1 vccd1 vccd1 y_r_3[13] sky130_fd_sc_hd__buf_2
Xoutput462 output462/A vssd1 vssd1 vccd1 vccd1 y_r_3[8] sky130_fd_sc_hd__buf_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput473 output473/A vssd1 vssd1 vccd1 vccd1 y_r_4[2] sky130_fd_sc_hd__buf_2
Xoutput484 output484/A vssd1 vssd1 vccd1 vccd1 y_r_5[12] sky130_fd_sc_hd__buf_2
XANTENNA__14789__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput495 _15617_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[7] sky130_fd_sc_hd__buf_2
XFILLER_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12894__A0 _13203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07989_ _11447_/B _08074_/C _11458_/A vssd1 vssd1 vccd1 vccd1 _07990_/B sky130_fd_sc_hd__mux2_1
XFILLER_170_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09728_ _09846_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _15718_/D sky130_fd_sc_hd__xnor2_1
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _09659_/A _09659_/B _09659_/C vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__and3_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A x_i_6[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12735_/C sky130_fd_sc_hd__xnor2_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07630__S _07632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ _11550_/A _11550_/B _11620_/X vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__a21o_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08617__A2 _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14029__A _14029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14340_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14359_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_169_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _15020_/Q vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_168_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ _15253_/Q _10502_/Y _10498_/B vssd1 vssd1 vccd1 vccd1 _10505_/B sky130_fd_sc_hd__a21o_1
X_11483_ _11483_/A _11483_/B vssd1 vssd1 vccd1 vccd1 _11564_/A sky130_fd_sc_hd__xnor2_1
X_14271_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14271_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input71_A x_i_4[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ _13222_/A _13222_/B vssd1 vssd1 vccd1 vccd1 _13240_/B sky130_fd_sc_hd__or2_1
X_10434_ _10434_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _14954_/D sky130_fd_sc_hd__xnor2_2
XFILLER_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10365_ _15133_/Q _15166_/Q vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__and2b_1
X_13153_ _13153_/A _13319_/A _13220_/A vssd1 vssd1 vccd1 vccd1 _13157_/A sky130_fd_sc_hd__and3_1
XFILLER_152_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10292__A _15153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ _12451_/B _12105_/B vssd1 vssd1 vccd1 vccd1 _12104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _13177_/A _13176_/A vssd1 vssd1 vccd1 vccd1 _13175_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10296_ _15152_/Q _10296_/B vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__nand2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14699__A _14701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12035_ _12038_/A _12122_/A _12055_/A vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__and3_1
XFILLER_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output325_A output325/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_890 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13986_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15725_ _15725_/CLK _15725_/D _14801_/Y vssd1 vssd1 vccd1 vccd1 _15725_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _12937_/A _12937_/B vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15656_ _15689_/CLK _15656_/D _14729_/Y vssd1 vssd1 vccd1 vccd1 _15656_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12868_ _12797_/B _12868_/B vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__and2b_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14607_/Y sky130_fd_sc_hd__inv_2
X_11819_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11821_/C sky130_fd_sc_hd__xnor2_1
XFILLER_187_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater642_A _11250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ _15784_/CLK _15587_/D _14656_/Y vssd1 vssd1 vccd1 vccd1 _15587_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12799_/A vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14538_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14538_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14469_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14469_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater907_A repeater908/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_938 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_908 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ _08961_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _15195_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07912_ _13591_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__and2_1
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14402__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ _15469_/Q _15453_/Q vssd1 vssd1 vccd1 vccd1 _08892_/X sky130_fd_sc_hd__and2b_1
XFILLER_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater910 input203/X vssd1 vssd1 vccd1 vccd1 _07864_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater921 input187/X vssd1 vssd1 vccd1 vccd1 _07702_/A1 sky130_fd_sc_hd__clkbuf_2
X_07843_ _07843_/A vssd1 vssd1 vccd1 vccd1 _15346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater932 input170/X vssd1 vssd1 vccd1 vccd1 _07834_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater943 input158/X vssd1 vssd1 vccd1 vccd1 _07761_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater954 input142/X vssd1 vssd1 vccd1 vccd1 _07890_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater965 input127/X vssd1 vssd1 vccd1 vccd1 _07400_/A1 sky130_fd_sc_hd__clkbuf_2
X_07774_ _07774_/A vssd1 vssd1 vccd1 vccd1 _15380_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater976 input116/X vssd1 vssd1 vccd1 vccd1 _07392_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _15532_/Q _15516_/Q _09512_/X vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12857__A _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _15532_/Q _15516_/Q vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__and2b_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11480__B _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09377_/B sky130_fd_sc_hd__and2_1
XFILLER_71_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_740 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ _08280_/Y _08342_/A vssd1 vssd1 vccd1 vccd1 _08326_/X sky130_fd_sc_hd__and2b_1
XFILLER_71_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ _08257_/A _08257_/B vssd1 vssd1 vccd1 vccd1 _08281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_166_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_180_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ _08190_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__xor2_1
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _10839_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _15802_/D sky130_fd_sc_hd__xnor2_1
XFILLER_133_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput270 output270/A vssd1 vssd1 vccd1 vccd1 y_i_0[3] sky130_fd_sc_hd__buf_2
Xoutput281 output281/A vssd1 vssd1 vccd1 vccd1 y_i_1[13] sky130_fd_sc_hd__buf_2
XFILLER_160_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput292 output292/A vssd1 vssd1 vccd1 vccd1 y_i_1[8] sky130_fd_sc_hd__buf_2
X_10081_ _10079_/X _10087_/A vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14312__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__A1 _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09406__A _15509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_646 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13840_ _13840_/A _13842_/B vssd1 vssd1 vccd1 vccd1 _15669_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input223_A x_r_5[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08299__B1 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13771_ _13783_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13772_/C sky130_fd_sc_hd__xor2_1
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _10982_/B _10982_/C _10982_/A vssd1 vssd1 vccd1 vccd1 _10984_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15510_ _15525_/CLK _15510_/D _14574_/Y vssd1 vssd1 vccd1 vccd1 _15510_/Q sky130_fd_sc_hd__dfrtp_1
X_12722_ _12723_/A _12726_/A _12723_/C vssd1 vssd1 vccd1 vccd1 _12836_/A sky130_fd_sc_hd__o21ai_1
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15441_ _15803_/CLK _15441_/D _14502_/Y vssd1 vssd1 vccd1 vccd1 _15441_/Q sky130_fd_sc_hd__dfrtp_2
X_12653_ _12653_/A _12726_/C vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11604_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15372_ _15724_/CLK _15372_/D _14428_/Y vssd1 vssd1 vccd1 vccd1 _15372_/Q sky130_fd_sc_hd__dfrtp_4
X_12584_ _12583_/A _12583_/B _12578_/B _12579_/Y _12580_/Y vssd1 vssd1 vccd1 vccd1
+ _12585_/B sky130_fd_sc_hd__o221ai_2
XFILLER_12_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_732 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11537_/C sky130_fd_sc_hd__xnor2_1
XFILLER_102_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14254_/Y sky130_fd_sc_hd__inv_2
X_11466_ _11466_/A _08196_/A vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__or2b_1
XFILLER_171_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output275_A output275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13205_ _13205_/A _13277_/B vssd1 vssd1 vccd1 vccd1 _13208_/A sky130_fd_sc_hd__xor2_4
XFILLER_125_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10417_ _10417_/A _10417_/B _10417_/C vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__and3_1
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14185_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14185_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11397_ _10202_/A _11396_/B _10202_/B vssd1 vssd1 vccd1 vccd1 _11398_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__12007__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_661 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13136_ _13138_/A _13138_/C vssd1 vssd1 vccd1 vccd1 _13137_/B sky130_fd_sc_hd__or2_1
X_10348_ _15130_/Q _15163_/Q vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output442_A output442/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13138_/A _13066_/Y vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__nor2b_1
X_10279_ _10279_/A _10279_/B _11424_/A vssd1 vssd1 vccd1 vccd1 _10281_/A sky130_fd_sc_hd__and3_1
XANTENNA__14222__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12018_ _12018_/A _12454_/B vssd1 vssd1 vccd1 vccd1 _12223_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13969_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12677__A _13431_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15708_ _15708_/CLK _15708_/D _14784_/Y vssd1 vssd1 vccd1 vccd1 _15708_/Q sky130_fd_sc_hd__dfrtp_1
X_07490_ _15519_/Q _07490_/A1 _07538_/S vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15639_ _15705_/CLK _15639_/D _14711_/Y vssd1 vssd1 vccd1 vccd1 _15639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09160_ _09639_/A _09160_/B vssd1 vssd1 vccd1 vccd1 _15288_/D sky130_fd_sc_hd__xnor2_1
X_08111_ _08305_/A vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__inv_2
XFILLER_148_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_771 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09091_ _09233_/A _09091_/B vssd1 vssd1 vccd1 vccd1 _15223_/D sky130_fd_sc_hd__xor2_1
XFILLER_174_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ _08060_/A _08060_/B _08041_/Y vssd1 vssd1 vccd1 vccd1 _08045_/A sky130_fd_sc_hd__a21oi_1
XFILLER_135_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09993_/A _09993_/B _09993_/C vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__nor3_1
XFILLER_153_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _15464_/Q _15448_/Q _08943_/X vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14132__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07445__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08130__A _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _15466_/Q _15450_/Q vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__and2b_1
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater740 _15660_/Q vssd1 vssd1 vccd1 vccd1 output311/A sky130_fd_sc_hd__buf_2
XANTENNA__13971__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater751 repeater752/X vssd1 vssd1 vccd1 vccd1 output292/A sky130_fd_sc_hd__buf_4
X_07826_ _15354_/Q input174/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07827_/A sky130_fd_sc_hd__mux2_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater762 _15640_/Q vssd1 vssd1 vccd1 vccd1 output520/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater773 _15625_/Q vssd1 vssd1 vccd1 vccd1 output487/A sky130_fd_sc_hd__clkbuf_2
Xrepeater784 _15608_/Q vssd1 vssd1 vccd1 vccd1 output452/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater795 _15594_/Q vssd1 vssd1 vccd1 vccd1 output447/A sky130_fd_sc_hd__clkbuf_2
X_07757_ _15388_/Q _07757_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08784__B _15323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11491__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ _07688_/A vssd1 vssd1 vccd1 vccd1 _15422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09427_ _15530_/Q _15514_/Q vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _09357_/Y _15383_/Q _09356_/B vssd1 vssd1 vccd1 vccd1 _09359_/B sky130_fd_sc_hd__a21o_1
XFILLER_12_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08309_ _08310_/A _08310_/B _08287_/X _08289_/X vssd1 vssd1 vccd1 vccd1 _08309_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14952__D _14952_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09289_ _09359_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _15122_/D sky130_fd_sc_hd__xor2_1
XFILLER_139_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14307__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ _11319_/B _11319_/C _11319_/A vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11251_ _11251_/A _11251_/B _11251_/C vssd1 vssd1 vccd1 vccd1 _11253_/A sky130_fd_sc_hd__and3_1
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input173_A x_r_2[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__nand2_2
XFILLER_84_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11182_ _11181_/A _11181_/C _11363_/A vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15783__D _15783_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11666__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _10125_/Y _10129_/B _10127_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__o21ai_1
XFILLER_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14042__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A _15297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14941_ _15732_/CLK _14941_/D _13972_/Y vssd1 vssd1 vccd1 vccd1 _14941_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_input34_A x_i_1[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _15212_/Q _15113_/Q vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__xor2_2
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13823_ _14975_/Q _13824_/B vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ _13741_/A _13741_/B _14980_/Q vssd1 vssd1 vccd1 vccd1 _13754_/Y sky130_fd_sc_hd__o21ai_1
X_10966_ _10966_/A _10966_/B _10966_/C vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__and3_1
XFILLER_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12705_ _12636_/A _12636_/B _12635_/A vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__a21oi_1
XFILLER_204_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ _14975_/Q vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__inv_2
X_10897_ _10897_/A _10902_/A vssd1 vssd1 vccd1 vccd1 _10897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15424_ _15438_/CLK _15424_/D _14484_/Y vssd1 vssd1 vccd1 vccd1 _15424_/Q sky130_fd_sc_hd__dfrtp_4
X_12636_ _12636_/A _12636_/B vssd1 vssd1 vccd1 vccd1 _12643_/A sky130_fd_sc_hd__xor2_1
XFILLER_15_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output392_A _15698_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _15722_/CLK _15355_/D _14410_/Y vssd1 vssd1 vccd1 vccd1 _15355_/Q sky130_fd_sc_hd__dfrtp_1
X_12567_ _12567_/A vssd1 vssd1 vccd1 vccd1 _12567_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14217__A _14218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13121__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14306_/Y sky130_fd_sc_hd__inv_2
X_11518_ _11588_/A _11588_/B vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__xor2_1
XFILLER_172_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15286_ _15592_/CLK _15286_/D _14337_/Y vssd1 vssd1 vccd1 vccd1 _15286_/Q sky130_fd_sc_hd__dfrtp_1
X_12498_ _12498_/A _12498_/B vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14237_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14237_/Y sky130_fd_sc_hd__inv_2
X_11449_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__xnor2_1
XFILLER_171_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater605_A _10753_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14168_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08869__B _15449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13025_/A _13025_/B _13036_/B _13041_/A vssd1 vssd1 vccd1 vccd1 _13120_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14099_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14118_/A sky130_fd_sc_hd__buf_12
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater974_A repeater975/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14887__A _14889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08660_ _12650_/B _08660_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07611_ _07611_/A vssd1 vssd1 vccd1 vccd1 _15460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08591_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08591_/X sky130_fd_sc_hd__or2_1
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07542_ _07542_/A vssd1 vssd1 vccd1 vccd1 _15494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ _15527_/Q _07473_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07474_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09212_ _09212_/A vssd1 vssd1 vccd1 vccd1 _09680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12854__B _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ _15542_/Q _15562_/Q vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__or2b_1
XFILLER_175_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__A _15273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14127__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13031__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09074_ _15495_/Q _15479_/Q vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__and2_1
XFILLER_190_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ _08025_/A _08025_/B _08025_/C vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or3_1
XANTENNA__13966__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08779__B _15322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A1 _07410_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09976_ _09880_/A _09975_/B _09880_/B vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__a21boi_1
XFILLER_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08927_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _15215_/D sky130_fd_sc_hd__nor2_1
XFILLER_190_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14797__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _15464_/Q _15448_/Q vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__xnor2_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater570 _11131_/X vssd1 vssd1 vccd1 vccd1 repeater570/X sky130_fd_sc_hd__buf_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater581 _11329_/Y vssd1 vssd1 vccd1 vccd1 repeater581/X sky130_fd_sc_hd__buf_2
XFILLER_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _07809_/A vssd1 vssd1 vccd1 vccd1 _15363_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14947__D _14947_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater592 _11061_/Y vssd1 vssd1 vccd1 vccd1 output276/A sky130_fd_sc_hd__clkbuf_2
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08789_ _15340_/Q _15324_/Q vssd1 vssd1 vccd1 vccd1 _13890_/A sky130_fd_sc_hd__xnor2_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _14909_/D sky130_fd_sc_hd__xor2_2
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07477__A1 _07477_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _10751_/A _10751_/B vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__nand2_4
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08019__B _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _13470_/A _13470_/B _13470_/C vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__and3_1
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10682_ _10679_/A _10999_/A _10679_/B _10681_/X vssd1 vssd1 vccd1 vccd1 _10685_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_90_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15778__D _15778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12421_ _12596_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12594_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14037__A _14037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15140_ _15406_/CLK _15140_/D _14183_/Y vssd1 vssd1 vccd1 vccd1 _15140_/Q sky130_fd_sc_hd__dfrtp_1
X_12352_ _14939_/Q vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__inv_2
XFILLER_5_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08035__A _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _11303_/A _11303_/B _11303_/C vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__and3_1
XFILLER_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15071_ _15352_/CLK _15071_/D _14110_/Y vssd1 vssd1 vccd1 vccd1 _15071_/Q sky130_fd_sc_hd__dfrtp_1
X_12283_ _12312_/S _12246_/X _12247_/B vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__o21ai_1
XFILLER_142_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12780__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08729__A1 _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14022_/Y sky130_fd_sc_hd__inv_2
X_11234_ _15756_/Q _15034_/Q vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__xor2_4
XFILLER_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11165_ _11163_/Y _11165_/B vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__and2b_1
XFILLER_171_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _15139_/Q _15304_/Q vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__nand2_1
X_11096_ _14935_/Q _15001_/Q _11095_/B vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__a21oi_1
XFILLER_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15018__D _15018_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ _15220_/CLK _14924_/D _13954_/Y vssd1 vssd1 vccd1 vccd1 _14924_/Q sky130_fd_sc_hd__dfrtp_1
X_10047_ _15209_/Q _15110_/Q vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__nand2_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14500__A _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14855_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output405_A output405/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _13806_/A _13806_/B vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14786_ _14787_/A vssd1 vssd1 vccd1 vccd1 _14786_/Y sky130_fd_sc_hd__inv_2
X_11998_ _11999_/A _11999_/B vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _13295_/B _13737_/B vssd1 vssd1 vccd1 vccd1 _13744_/B sky130_fd_sc_hd__and2b_1
XFILLER_188_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10949_ _14968_/Q _14902_/Q vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__xor2_4
XFILLER_43_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater555_A repeater556/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clkbuf_opt_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _15687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13668_ _13677_/C _13668_/B vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12674__B _12970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15407_ _15808_/CLK _15407_/D _14466_/Y vssd1 vssd1 vccd1 vccd1 _15407_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _14953_/Q _12620_/B vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__and2_1
XFILLER_192_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater722_A _15693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13599_ _15368_/Q _15352_/Q _13598_/X vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ _15722_/CLK _15338_/D _14392_/Y vssd1 vssd1 vccd1 vccd1 _15338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_583 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07640__A1 _07640_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ _15561_/CLK _15269_/D _14319_/Y vssd1 vssd1 vccd1 vccd1 _15269_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09830_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09832_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09761_ _09760_/A _09760_/B _09861_/A vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__a21oi_1
XFILLER_140_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09145__A1 _15561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ _08748_/B _08710_/X _08748_/A vssd1 vssd1 vccd1 vccd1 _08712_/Y sky130_fd_sc_hd__a21oi_1
X_09692_ _09690_/Y _09692_/B vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__and2b_1
XANTENNA__14410__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _12654_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13026__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12482__B_N _12213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _08598_/A _08596_/A _08621_/A vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__or3_1
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07525_/A vssd1 vssd1 vccd1 vccd1 _15502_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07459__A1 _07459_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07959__A _15251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_354 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07456_ _07456_/A vssd1 vssd1 vccd1 vccd1 _15536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07387_ _07387_/A vssd1 vssd1 vccd1 vccd1 _15574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ _15505_/Q _15489_/Q vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__and2_1
XFILLER_157_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09057_ _09056_/A _09056_/B _13628_/A vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__o21a_1
XFILLER_203_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08008_ _11447_/B _11458_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__and3_1
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12105__A _12451_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _09958_/A _09958_/B _10003_/A vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__a21oi_1
XFILLER_106_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _12970_/A _12970_/B vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__xnor2_4
XFILLER_57_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input136_A x_r_0[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14320__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ _11921_/A _11921_/B vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11663__B _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14640_/Y sky130_fd_sc_hd__inv_2
X_11852_ _11852_/A _11852_/B vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__or2_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _15724_/Q _15790_/Q vssd1 vssd1 vccd1 vccd1 _10803_/Y sky130_fd_sc_hd__nand2_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14571_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14571_/Y sky130_fd_sc_hd__inv_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11783_/A _11783_/B _12391_/B vssd1 vssd1 vccd1 vccd1 _11787_/B sky130_fd_sc_hd__or3b_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15694_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13522_ _13522_/A vssd1 vssd1 vccd1 vccd1 _13522_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10734_ _15713_/Q _15779_/Q vssd1 vssd1 vccd1 vccd1 _10734_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__A1 _07870_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ _13770_/B _13770_/A vssd1 vssd1 vccd1 vccd1 _13453_/X sky130_fd_sc_hd__or2b_1
XFILLER_201_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10665_ _15275_/Q _15176_/Q vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12404_ _12391_/A _12391_/B _12403_/X vssd1 vssd1 vccd1 vccd1 _12406_/C sky130_fd_sc_hd__o21a_1
XFILLER_142_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _13384_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _13385_/B sky130_fd_sc_hd__and2_1
XFILLER_12_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10596_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _14991_/D sky130_fd_sc_hd__xnor2_1
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15123_ _15406_/CLK _15123_/D _14165_/Y vssd1 vssd1 vccd1 vccd1 _15123_/Q sky130_fd_sc_hd__dfrtp_1
X_12335_ _12335_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12335_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07622__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_705 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07808__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15054_ _15352_/CLK _15054_/D _14092_/Y vssd1 vssd1 vccd1 vccd1 _15054_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ _15738_/Q _12564_/B vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__xnor2_1
XFILLER_99_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output355_A output355/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14005_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14005_/Y sky130_fd_sc_hd__inv_2
X_11217_ _11216_/A _11216_/B _11375_/A vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__a21o_1
X_12197_ _12198_/B _12197_/B vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12015__A _12439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11148_ _11248_/A _14987_/Q _11353_/B vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__a21o_1
XANTENNA_output522_A output522/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_635 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _11077_/X _11085_/A vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14230__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput170 x_r_2[1] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__clkbuf_1
Xinput181 x_r_3[11] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_hd__clkbuf_2
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07543__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput192 x_r_3[7] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07689__A1 _07689_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ _15400_/CLK _14907_/D _13936_/Y vssd1 vssd1 vccd1 vccd1 _14907_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_repeater672_A _14675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ _14841_/A vssd1 vssd1 vccd1 vccd1 _14838_/Y sky130_fd_sc_hd__inv_2
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14769_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14769_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_43_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _15170_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08290_ _11797_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__or2_1
XFILLER_60_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_870 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14405__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A_N _15446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09813_ _09620_/A _09812_/B _09620_/B vssd1 vssd1 vccd1 vccd1 _15168_/D sky130_fd_sc_hd__a21boi_1
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07961__B _15251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _09744_/A _09744_/B _09857_/A vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__and3_1
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14140__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07453__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09675_ _09675_/A _09675_/B _09675_/C vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__and3_1
XFILLER_27_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08617_/X _08622_/Y _08722_/B _08724_/B _08742_/B vssd1 vssd1 vccd1 vccd1
+ _08626_/X sky130_fd_sc_hd__o311a_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08557_ _08566_/A _08566_/B vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15392_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08792__B _08792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07508_ _15510_/Q input26/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08488_ _12780_/A _08478_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08488_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_966 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07852__A1 input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ _15544_/Q _07439_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07440_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12189__B1 _12312_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10450_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _14893_/D sky130_fd_sc_hd__xor2_1
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ _09245_/A _09113_/B vssd1 vssd1 vccd1 vccd1 _15227_/D sky130_fd_sc_hd__xor2_1
XFILLER_184_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14960__D _14960_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A1 _07604_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ _15086_/Q _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10383_/C sky130_fd_sc_hd__a21o_1
XFILLER_191_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14315__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ _12181_/A _12120_/B vssd1 vssd1 vccd1 vccd1 _12122_/B sky130_fd_sc_hd__and2_1
XANTENNA__07628__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ _12119_/B _12051_/B vssd1 vssd1 vccd1 vccd1 _12053_/C sky130_fd_sc_hd__or2_1
XFILLER_172_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input253_A x_r_7[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08032__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _11002_/A vssd1 vssd1 vccd1 vccd1 _15014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15810_ _15810_/A vssd1 vssd1 vccd1 vccd1 _15810_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14050__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _15741_/CLK _15741_/D _14818_/Y vssd1 vssd1 vccd1 vccd1 _15741_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_891 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _13390_/A _13319_/A _12953_/C vssd1 vssd1 vccd1 vccd1 _13116_/B sky130_fd_sc_hd__and3_1
XANTENNA__12664__A1 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11904_/A _11904_/B vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _15707_/CLK _15672_/D _14746_/Y vssd1 vssd1 vccd1 vccd1 _15672_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12824_/S _12921_/A _13201_/A _12714_/B _13012_/A vssd1 vssd1 vccd1 vccd1
+ _12884_/X sky130_fd_sc_hd__o2111a_1
XFILLER_18_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__A _15365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14623_/Y sky130_fd_sc_hd__inv_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11835_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__nor2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15279_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14554_/Y sky130_fd_sc_hd__inv_2
X_11766_ _11766_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10978__A1 _15271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13505_ _13505_/A _13505_/B vssd1 vssd1 vccd1 vccd1 _13506_/S sky130_fd_sc_hd__nand2_1
X_10717_ _10717_/A _11016_/A vssd1 vssd1 vccd1 vccd1 _15052_/D sky130_fd_sc_hd__xnor2_4
X_14485_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__inv_2
X_11697_ _11928_/A _12088_/A _11697_/C vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__and3_1
XFILLER_158_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13436_ _13455_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__xor2_1
X_10648_ _10642_/A _10644_/B _10642_/B vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__a21boi_4
XFILLER_42_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output472_A output472/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12952__B _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11849__A _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13367_ _13425_/B _13367_/B vssd1 vssd1 vccd1 vccd1 _13369_/C sky130_fd_sc_hd__nand2_1
XANTENNA__14225__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ _10579_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _15034_/D sky130_fd_sc_hd__nor2_1
XFILLER_155_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15367_/CLK _15106_/D _14147_/Y vssd1 vssd1 vccd1 vccd1 _15106_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__07538__S _07538_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ _12319_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_895 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08223__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13298_ _13352_/A _13298_/B vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__nand2_1
X_15037_ _15525_/CLK _15037_/D _14074_/Y vssd1 vssd1 vccd1 vccd1 _15037_/Q sky130_fd_sc_hd__dfrtp_1
X_12249_ _12190_/A _12247_/Y _12246_/X _12245_/Y vssd1 vssd1 vccd1 vccd1 _12250_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_64_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater887_A input237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _07790_/A vssd1 vssd1 vccd1 vccd1 _15372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15206__D _15206_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ _09459_/A _09459_/B _09518_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08411_ _08411_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08429_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09391_ _09390_/A _09390_/C _09390_/B vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__a21oi_1
XFILLER_196_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _15221_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_205_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08342_ _08342_/A _08280_/Y vssd1 vssd1 vccd1 vccd1 _08342_/X sky130_fd_sc_hd__or2b_1
XFILLER_205_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_944 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08273_ _08273_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _08321_/B sky130_fd_sc_hd__xnor2_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07834__A1 _07834_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_969 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11759__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07598__A0 _15466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14135__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__A _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput430 output430/A vssd1 vssd1 vccd1 vccd1 y_r_2[0] sky130_fd_sc_hd__buf_2
Xoutput441 output441/A vssd1 vssd1 vccd1 vccd1 y_r_2[4] sky130_fd_sc_hd__buf_2
XFILLER_195_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13974__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput452 output452/A vssd1 vssd1 vccd1 vccd1 y_r_3[14] sky130_fd_sc_hd__buf_2
XFILLER_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_888 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput463 output463/A vssd1 vssd1 vccd1 vccd1 y_r_3[9] sky130_fd_sc_hd__buf_2
Xoutput474 _11256_/X vssd1 vssd1 vccd1 vccd1 y_r_4[3] sky130_fd_sc_hd__buf_2
Xoutput485 _15623_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[13] sky130_fd_sc_hd__buf_2
Xoutput496 output496/A vssd1 vssd1 vccd1 vccd1 y_r_5[8] sky130_fd_sc_hd__buf_2
XFILLER_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13185__S _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07988_ _11584_/A vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__inv_2
XFILLER_41_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _09719_/Y _09723_/B _09721_/B vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__o21ai_2
XFILLER_41_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ _15570_/Q _15550_/Q vssd1 vssd1 vccd1 vccd1 _09659_/C sky130_fd_sc_hd__or2b_1
XFILLER_103_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07522__A0 _15503_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _08603_/X _08606_/X _08732_/A vssd1 vssd1 vccd1 vccd1 _08609_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_747 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09589_ _09589_/A _09597_/A vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__nand2_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11620_ _11549_/B _11620_/B vssd1 vssd1 vccd1 vccd1 _11620_/X sky130_fd_sc_hd__and2b_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09814__A2 _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ _12247_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__nand2_1
XFILLER_211_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10502_ _15286_/Q vssd1 vssd1 vccd1 vccd1 _10502_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14270_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14270_/Y sky130_fd_sc_hd__inv_2
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11483_/B sky130_fd_sc_hd__xor2_1
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13221_ _13221_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13240_/A sky130_fd_sc_hd__or2_1
XANTENNA__11669__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ _10432_/A _10432_/B _10093_/B vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07589__A0 _15470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14045__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13152_ _13330_/A _13152_/B vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__nand2_1
XANTENNA_input64_A x_i_3[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10364_ _15132_/Q _15165_/Q vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _12096_/B _12096_/C _15735_/Q vssd1 vssd1 vccd1 vccd1 _12156_/B sky130_fd_sc_hd__a21bo_1
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13083_ _13083_/A _13083_/B vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__xnor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10295_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _15776_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__08978__A _15349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _12178_/A vssd1 vssd1 vccd1 vccd1 _12038_/A sky130_fd_sc_hd__inv_2
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13985_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1019 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output318_A output318/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15724_ _15724_/CLK _15724_/D _14800_/Y vssd1 vssd1 vccd1 vccd1 _15724_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12936_ _12991_/A _12991_/B vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__A _15441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _15690_/CLK _15655_/D _14728_/Y vssd1 vssd1 vccd1 vccd1 _15655_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12867_ _12867_/A _12867_/B vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__xnor2_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _11901_/A _11818_/B vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__and2_1
XFILLER_18_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14606_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__inv_2
X_15586_ _15784_/CLK _15586_/D _14655_/Y vssd1 vssd1 vccd1 vccd1 _15586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__A _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ _12798_/A _12798_/B vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__xor2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07816__A1 _07816_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14537_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14537_/Y sky130_fd_sc_hd__inv_2
X_11749_ _11749_/A _11749_/B _11749_/C vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__and3_1
XFILLER_187_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater635_A repeater636/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14468_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14468_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15696__D _15696_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ _13419_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__xnor2_1
XFILLER_162_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater802_A _15588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14399_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14399_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ _08959_/A _08959_/C _08959_/B vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_5_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _15573_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08888__A _15470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07911_ _15365_/Q _15349_/Q vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__or2_1
XFILLER_151_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08891_ _08891_/A vssd1 vssd1 vccd1 vccd1 _08957_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater900 input220/X vssd1 vssd1 vccd1 vccd1 _07732_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater911 input202/X vssd1 vssd1 vccd1 vccd1 _07866_/A1 sky130_fd_sc_hd__buf_4
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07842_ _15346_/Q _07842_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07843_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater922 repeater923/X vssd1 vssd1 vccd1 vccd1 _07704_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__12203__A _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater933 input17/X vssd1 vssd1 vccd1 vccd1 _07624_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater944 input157/X vssd1 vssd1 vccd1 vccd1 _07763_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater955 input141/X vssd1 vssd1 vccd1 vccd1 _07892_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater966 input125/X vssd1 vssd1 vccd1 vccd1 _07404_/A1 sky130_fd_sc_hd__buf_4
X_07773_ _15380_/Q _07773_/A1 _07791_/S vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__mux2_1
Xrepeater977 input115/X vssd1 vssd1 vccd1 vccd1 _07412_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_186_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_861 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09512_ _15532_/Q _15516_/Q _09511_/B vssd1 vssd1 vccd1 vccd1 _09512_/X sky130_fd_sc_hd__o21a_1
XFILLER_209_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07504__A0 _15512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12857__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _09441_/Y _09443_/B vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__nand2b_2
XFILLER_24_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__C _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _15143_/D sky130_fd_sc_hd__xor2_1
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08325_ _08325_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__xor2_1
XFILLER_127_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13969__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ _08307_/A vssd1 vssd1 vccd1 vccd1 _08281_/A sky130_fd_sc_hd__inv_2
XFILLER_193_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09068__B_N _15494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08187_ _12204_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08190_/B sky130_fd_sc_hd__xnor2_1
XFILLER_134_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_81_clk_A _14904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput260 _15810_/A vssd1 vssd1 vccd1 vccd1 y_i_0[0] sky130_fd_sc_hd__buf_2
Xoutput271 output271/A vssd1 vssd1 vccd1 vccd1 y_i_0[4] sky130_fd_sc_hd__buf_2
XANTENNA__13323__A_N _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput282 output282/A vssd1 vssd1 vccd1 vccd1 y_i_1[14] sky130_fd_sc_hd__buf_2
XFILLER_160_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput293 output293/A vssd1 vssd1 vccd1 vccd1 y_i_1[9] sky130_fd_sc_hd__buf_2
XFILLER_47_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10079_/A _10079_/B _10428_/A vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_96_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__A2 _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13209__A _13722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08905__B_N _15456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_774 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12113__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11952__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08299__A1 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13770_ _13770_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13783_/A sky130_fd_sc_hd__nor2_1
XANTENNA_input216_A x_r_5[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08299__B2 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _10982_/A _10982_/B _10982_/C vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__and3_1
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12721_ _12812_/A _12721_/B vssd1 vssd1 vccd1 vccd1 _12723_/C sky130_fd_sc_hd__xnor2_1
XFILLER_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09422__A _15529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ _15699_/CLK _15440_/D _14500_/Y vssd1 vssd1 vccd1 vccd1 _15440_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _12652_/A _12652_/B vssd1 vssd1 vccd1 vccd1 _12726_/C sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__xnor2_1
X_15371_ _15617_/CLK _15371_/D _14427_/Y vssd1 vssd1 vccd1 vccd1 _15371_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13595__A2 _15351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11534_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__xor2_1
XFILLER_128_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_935 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14253_/Y sky130_fd_sc_hd__inv_2
X_11465_ _08269_/A _08269_/B _11464_/X vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_49_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ _13197_/B _13090_/B _13093_/B _13203_/X vssd1 vssd1 vccd1 vccd1 _13277_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10416_ _15111_/Q _15210_/Q vssd1 vssd1 vccd1 vccd1 _10417_/C sky130_fd_sc_hd__or2b_1
X_14184_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14184_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _11396_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _15729_/D sky130_fd_sc_hd__xnor2_1
XFILLER_48_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output268_A _11020_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ _12981_/A _13547_/A _12982_/Y _13066_/Y vssd1 vssd1 vccd1 vccd1 _13138_/C
+ sky130_fd_sc_hd__o211a_1
X_10347_ _10347_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__nand2_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14503__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07816__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13066_ _15764_/Q _13066_/B vssd1 vssd1 vccd1 vccd1 _13066_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08501__A _15792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _15083_/Q _15248_/Q vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__xor2_4
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output435_A output435/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _11940_/A _11940_/B _11951_/Y _11952_/Y vssd1 vssd1 vccd1 vccd1 _12018_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_107_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13968_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13968_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07551__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15707_ _15707_/CLK _15707_/D _14783_/Y vssd1 vssd1 vccd1 vccd1 _15707_/Q sky130_fd_sc_hd__dfrtp_1
X_12919_ _15762_/Q _13545_/B vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__and2_1
XFILLER_179_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13899_ _13899_/A _13901_/B vssd1 vssd1 vccd1 vccd1 _15063_/D sky130_fd_sc_hd__nor2_1
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15638_ _15648_/CLK _15638_/D _14710_/Y vssd1 vssd1 vccd1 vccd1 _15638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _15569_/CLK _15569_/D _14636_/Y vssd1 vssd1 vccd1 vccd1 _15569_/Q sky130_fd_sc_hd__dfrtp_1
X_08110_ _08304_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08305_/A sky130_fd_sc_hd__nor2_1
XFILLER_202_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ _15497_/Q _15481_/Q _09089_/X vssd1 vssd1 vccd1 vccd1 _09091_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08041_ _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_703 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10941__A _10941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _15195_/Q _15228_/Q vssd1 vssd1 vccd1 vccd1 _09993_/C sky130_fd_sc_hd__and2_1
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14413__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07726__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08943_ _15464_/Q _15448_/Q _08942_/B vssd1 vssd1 vccd1 vccd1 _08943_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15666_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_9_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ _08872_/Y _08874_/B vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__nand2b_2
XFILLER_28_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08130__B _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater730 _15678_/Q vssd1 vssd1 vccd1 vccd1 output354/A sky130_fd_sc_hd__clkbuf_2
Xrepeater741 _15659_/Q vssd1 vssd1 vccd1 vccd1 output284/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _07825_/A vssd1 vssd1 vccd1 vccd1 _15355_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater752 _15651_/Q vssd1 vssd1 vccd1 vccd1 repeater752/X sky130_fd_sc_hd__buf_2
Xrepeater763 _15639_/Q vssd1 vssd1 vccd1 vccd1 output519/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater774 _15624_/Q vssd1 vssd1 vccd1 vccd1 output486/A sky130_fd_sc_hd__clkbuf_2
Xrepeater785 _15607_/Q vssd1 vssd1 vccd1 vccd1 output451/A sky130_fd_sc_hd__clkbuf_2
X_07756_ _07756_/A vssd1 vssd1 vccd1 vccd1 _15389_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater796 repeater797/X vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07461__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _15422_/Q input194/X _07687_/S vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _09504_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _15271_/D sky130_fd_sc_hd__xor2_1
XFILLER_125_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09357_ _15399_/Q vssd1 vssd1 vccd1 vccd1 _09357_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08308_ _08308_/A vssd1 vssd1 vccd1 vccd1 _08310_/B sky130_fd_sc_hd__inv_2
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ _09284_/A _09283_/B _09283_/A vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__o21ba_1
XFILLER_166_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08239_ _08239_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08254_/A sky130_fd_sc_hd__nand2_1
XFILLER_154_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13211__B _13563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12108__A _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ _07969_/A _11248_/Y _11251_/C vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__o21a_2
XFILLER_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _15072_/Q _15237_/Q vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__nand2_1
XFILLER_192_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11181_ _11181_/A _11363_/A _11181_/C vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__and3_1
XFILLER_107_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14323__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input166_A x_r_2[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07636__S _07640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11666__B _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14940_ _15729_/CLK _14940_/D _13971_/Y vssd1 vssd1 vccd1 vccd1 _14940_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_85_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10063_ _10060_/A _10417_/A _10060_/B _10062_/X vssd1 vssd1 vccd1 vccd1 _10066_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A x_i_1[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14871_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_978 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13822_ _13822_/A _13822_/B vssd1 vssd1 vccd1 vccd1 _15665_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13753_ _13753_/A vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10965_ _07960_/A _10963_/Y _10966_/C vssd1 vssd1 vccd1 vccd1 _15005_/D sky130_fd_sc_hd__o21a_1
X_12704_ _12704_/A _12704_/B vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__and2_1
XFILLER_43_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13684_ _13684_/A _13822_/A vssd1 vssd1 vccd1 vccd1 _15697_/D sky130_fd_sc_hd__xor2_1
X_10896_ _10895_/A _10895_/C _11115_/A vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_599 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15423_ _15439_/CLK _15423_/D _14483_/Y vssd1 vssd1 vccd1 vccd1 _15423_/Q sky130_fd_sc_hd__dfrtp_1
X_12635_ _12635_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15354_ _15354_/CLK _15354_/D _14409_/Y vssd1 vssd1 vccd1 vccd1 _15354_/Q sky130_fd_sc_hd__dfrtp_2
X_12566_ _12566_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _15623_/D sky130_fd_sc_hd__xnor2_1
XFILLER_141_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output385_A output385/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _11517_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11588_/B sky130_fd_sc_hd__xnor2_1
X_14305_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14305_/Y sky130_fd_sc_hd__inv_2
X_15285_ _15592_/CLK _15285_/D _14336_/Y vssd1 vssd1 vccd1 vccd1 _15285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12497_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__or2_1
XFILLER_156_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14236_/Y sky130_fd_sc_hd__inv_2
X_11448_ _08010_/Y _11584_/A _11447_/X vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11857__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14167_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14233__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _11379_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__xor2_2
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13118_/B vssd1 vssd1 vccd1 vccd1 _13144_/B sky130_fd_sc_hd__xor2_1
XFILLER_113_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14098_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14098_/Y sky130_fd_sc_hd__inv_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _12970_/A _12970_/B _13048_/X vssd1 vssd1 vccd1 vccd1 _13050_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12688__A _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater967_A repeater968/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08885__B _15452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _15460_/Q _07610_/A1 _07632_/S vssd1 vssd1 vccd1 vccd1 _07611_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08590_ _08631_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08713_/B sky130_fd_sc_hd__xor2_2
XFILLER_53_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_8
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07541_ _15494_/Q input106/X _07591_/S vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07472_ _07472_/A vssd1 vssd1 vccd1 vccd1 _15528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__or2_1
XFILLER_50_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14408__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ _15562_/Q _15542_/Q vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__or2b_1
XANTENNA__13312__A _13357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ _15494_/Q _15478_/Q _09072_/B vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__a21oi_2
XFILLER_194_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08024_ _08025_/B _08025_/C _08025_/A vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__o21a_1
XFILLER_107_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10671__A _15276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14143__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _14924_/D sky130_fd_sc_hd__xnor2_1
XFILLER_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13982__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _08925_/A _08925_/B _08973_/A vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__o21a_1
XFILLER_170_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _15203_/D sky130_fd_sc_hd__nor2_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater560 _11382_/X vssd1 vssd1 vccd1 vccd1 output434/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07808_ _15363_/Q _07808_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__mux2_1
Xrepeater571 repeater572/X vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__buf_4
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater582 _11277_/Y vssd1 vssd1 vccd1 vccd1 output479/A sky130_fd_sc_hd__clkbuf_2
X_08788_ _13888_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _15075_/D sky130_fd_sc_hd__xor2_1
Xrepeater593 _10763_/Y vssd1 vssd1 vccd1 vccd1 output412/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _07739_/A vssd1 vssd1 vccd1 vccd1 _15397_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10750_ _15716_/Q _15782_/Q vssd1 vssd1 vccd1 vccd1 _10751_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ _09414_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__or2_1
XFILLER_200_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14963__D _14963_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10681_ _15277_/Q _15178_/Q vssd1 vssd1 vccd1 vccd1 _10681_/X sky130_fd_sc_hd__and2_1
XFILLER_129_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14318__A _14319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12420_ _12420_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__or2_1
XFILLER_185_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _12351_/A _12573_/A vssd1 vssd1 vccd1 vccd1 _15593_/D sky130_fd_sc_hd__xnor2_1
XFILLER_5_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08035__B _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _14921_/Q _11021_/Y _11303_/C vssd1 vssd1 vccd1 vccd1 _11302_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15070_ _15352_/CLK _15070_/D _14109_/Y vssd1 vssd1 vccd1 vccd1 _15070_/Q sky130_fd_sc_hd__dfrtp_1
X_12282_ _12190_/A _12245_/Y _12246_/X _12312_/S vssd1 vssd1 vccd1 vccd1 _12284_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15794__D _15794_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _14029_/A vssd1 vssd1 vccd1 vccd1 _14021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08729__A2 _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _11233_/A vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14053__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1004 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ _15746_/Q _15024_/Q vssd1 vssd1 vccd1 vccd1 _11165_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ _15139_/Q _15304_/Q vssd1 vssd1 vccd1 vccd1 _10115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11095_/Y sky130_fd_sc_hd__nor2_2
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _15119_/CLK _14923_/D _13953_/Y vssd1 vssd1 vccd1 vccd1 _14923_/Q sky130_fd_sc_hd__dfrtp_1
X_10046_ _15209_/Q _15110_/Q vssd1 vssd1 vccd1 vccd1 _10046_/Y sky130_fd_sc_hd__nor2_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _14861_/A vssd1 vssd1 vccd1 vccd1 _14854_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _14986_/Q _13805_/B vssd1 vssd1 vccd1 vccd1 _13806_/B sky130_fd_sc_hd__xnor2_1
XFILLER_17_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output300_A output300/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ _11997_/A _11997_/B vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__xnor2_1
XFILLER_189_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14785_ _14787_/A vssd1 vssd1 vccd1 vccd1 _14785_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10948_ _10948_/A vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__clkbuf_1
X_13736_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13744_/A sky130_fd_sc_hd__xor2_1
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879_ _10877_/Y _10879_/B vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__and2b_1
X_13667_ _13677_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__nand2_2
XANTENNA__14228__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15406_/CLK _15406_/D _14465_/Y vssd1 vssd1 vccd1 vccd1 _15406_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ _12618_/A _12618_/B vssd1 vssd1 vccd1 vccd1 _15691_/D sky130_fd_sc_hd__xor2_1
XFILLER_157_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08226__A _12088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _15368_/Q _15352_/Q _13597_/B vssd1 vssd1 vccd1 vccd1 _13598_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12549_ _12549_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__nand2_1
X_15337_ _15763_/CLK _15337_/D _14391_/Y vssd1 vssd1 vccd1 vccd1 _15337_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_repeater715_A _15704_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A1 _15497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15268_ _15268_/CLK _15268_/D _14318_/Y vssd1 vssd1 vccd1 vccd1 _15268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11587__A _11898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14238_/A sky130_fd_sc_hd__buf_12
XFILLER_99_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15199_ _15472_/CLK _15199_/D _14246_/Y vssd1 vssd1 vccd1 vccd1 _15199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _09760_/A _09760_/B _09861_/A vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__and3_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08896__A _15470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__and2_1
XFILLER_67_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09145__A2 _15541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _15055_/Q _15088_/Q vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _08426_/A _08640_/X _08641_/X vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__a21oi_1
XFILLER_55_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1017 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13026__B _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _08573_/A _08573_/B _08615_/A vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__or3_2
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07524_ _15502_/Q _07524_/A1 _07532_/S vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_683 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ _15536_/Q _07455_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_839 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__A _15275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14138__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07386_ _15574_/Q _07386_/A1 _07432_/S vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08136__A _11467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _09125_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _15230_/D sky130_fd_sc_hd__xor2_1
XFILLER_202_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13977__A _13977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12881__A _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09056_ _09056_/A _09056_/B _13628_/A vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__nor3_1
XFILLER_194_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08007_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08025_/C sky130_fd_sc_hd__and2_1
XFILLER_190_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _09958_/A _09958_/B _10003_/A vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__and3_1
XFILLER_66_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ _08907_/X _08914_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__and2b_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09889_/A _09977_/A _09889_/C vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__and3_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13217__A _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11920_ _11920_/A _11920_/B vssd1 vssd1 vccd1 vccd1 _11921_/B sky130_fd_sc_hd__nand2_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input129_A x_i_7[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11852_/A _11852_/B vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__nand2_1
XFILLER_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10802_/A _11298_/A vssd1 vssd1 vccd1 vccd1 _10802_/X sky130_fd_sc_hd__xor2_4
XFILLER_14_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14580_/A vssd1 vssd1 vccd1 vccd1 _14570_/Y sky130_fd_sc_hd__inv_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11782_ _12403_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__xnor2_2
XFILLER_26_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08647__A1 _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10733_ _11257_/A _10733_/B vssd1 vssd1 vccd1 vccd1 _10733_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_25_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ _13416_/A _13506_/S _15052_/Q vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__a21bo_1
XFILLER_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14048__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13452_ _13452_/A _13579_/A vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__nand2_1
XANTENNA_input94_A x_i_5[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ _10988_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _15043_/D sky130_fd_sc_hd__xnor2_4
XFILLER_9_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12403_ _12403_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _12403_/X sky130_fd_sc_hd__or2_1
XFILLER_173_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_990 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ _13384_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _13385_/A sky130_fd_sc_hd__nor2_1
XFILLER_142_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ _10501_/A _10594_/B _10501_/B vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__12791__A _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12334_ _12335_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15122_ _15279_/CLK _15122_/D _14164_/Y vssd1 vssd1 vccd1 vccd1 _15122_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_717 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15053_ _15477_/CLK _15053_/D _14091_/Y vssd1 vssd1 vccd1 vccd1 _15053_/Q sky130_fd_sc_hd__dfrtp_2
X_12265_ _12484_/A _12265_/B vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__xor2_2
XFILLER_154_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _14017_/A vssd1 vssd1 vccd1 vccd1 _14004_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11216_ _11216_/A _11216_/B _11375_/A vssd1 vssd1 vccd1 vccd1 _11216_/X sky130_fd_sc_hd__and3_1
X_12196_ _12254_/A _12131_/Y _12133_/A _12195_/Y vssd1 vssd1 vccd1 vccd1 _12197_/B
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__07386__A1 _07386_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output348_A _15688_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11147_ _14987_/Q _11353_/B vssd1 vssd1 vccd1 vccd1 _11147_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14511__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ _11077_/A _11077_/B _11344_/A vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__a21o_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput160 x_r_1[7] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_6
XFILLER_37_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput171 x_r_2[2] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput182 x_r_3[12] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14906_ _15399_/CLK _14906_/D _13935_/Y vssd1 vssd1 vccd1 vccd1 _14906_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_37_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10029_ _10023_/A _10025_/B _10023_/B vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__a21boi_2
Xinput193 x_r_3[8] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_2
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14837_ _14841_/A vssd1 vssd1 vccd1 vccd1 _14837_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater665_A _14753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14768_ _14781_/A vssd1 vssd1 vccd1 vccd1 _14768_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15699__D _15699_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater832_A repeater833/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ _13725_/B _13719_/B vssd1 vssd1 vccd1 vccd1 _13836_/B sky130_fd_sc_hd__nand2_1
XFILLER_204_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10486__A _10486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14699_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14699_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_642 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _15167_/D sky130_fd_sc_hd__xnor2_1
XFILLER_114_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_783 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14421__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07734__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11764__B _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13037__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09675_/C sky130_fd_sc_hd__nand2_1
XFILLER_28_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__or2b_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__xnor2_2
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07507_ _07507_/A vssd1 vssd1 vccd1 vccd1 _15511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1006 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08487_ _08728_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1028 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07438_ _07438_/A vssd1 vssd1 vccd1 vccd1 _15545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_978 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12189__A1 _12254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09108_ _15501_/Q _15485_/Q _09107_/X vssd1 vssd1 vccd1 vccd1 _09113_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _09038_/A _09038_/B _13618_/A vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _12050_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11001_ _10999_/X _11003_/C vssd1 vssd1 vccd1 vccd1 _11002_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input246_A x_r_7[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14331__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07644__S _07644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_915 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740_ _15741_/CLK _15740_/D _14817_/Y vssd1 vssd1 vccd1 vccd1 _15740_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _13438_/A _13381_/B vssd1 vssd1 vccd1 vccd1 _12953_/C sky130_fd_sc_hd__xor2_1
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__nand2_2
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _15708_/CLK _15671_/D _14745_/Y vssd1 vssd1 vccd1 vccd1 _15671_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12830_/B _12883_/B vssd1 vssd1 vccd1 vccd1 _12902_/B sky130_fd_sc_hd__and2b_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14640_/A vssd1 vssd1 vccd1 vccd1 _14622_/Y sky130_fd_sc_hd__inv_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11855_/B sky130_fd_sc_hd__or2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11765_ _11806_/C _11587_/B _11898_/A vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__mux2_1
XFILLER_144_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14553_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14553_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10716_ _15283_/Q _15184_/Q vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__xnor2_4
X_13504_ _13352_/A _13417_/B _13417_/A vssd1 vssd1 vccd1 vccd1 _13504_/X sky130_fd_sc_hd__a21o_1
XFILLER_18_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11696_ _11906_/A _11696_/B vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__nor2_1
XFILLER_202_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14484_ _14494_/A vssd1 vssd1 vccd1 vccd1 _14484_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13377__B1 _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10647_ _10645_/Y _10647_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__and2b_2
XFILLER_158_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ _13435_/A _13435_/B vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14506__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13366_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13367_/B sky130_fd_sc_hd__or2_1
XFILLER_127_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ _10577_/A _10577_/B _10622_/A vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__a21oi_1
X_15105_ _15367_/CLK _15105_/D _14146_/Y vssd1 vssd1 vccd1 vccd1 _15105_/Q sky130_fd_sc_hd__dfrtp_1
X_12317_ _12502_/A _12317_/B vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__xnor2_2
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297_ _13297_/A vssd1 vssd1 vccd1 vccd1 _13298_/B sky130_fd_sc_hd__inv_2
XANTENNA__12026__A _12439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08223__B _08223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12248_ _12245_/Y _12246_/X _12247_/Y _12190_/A vssd1 vssd1 vccd1 vccd1 _12250_/A
+ sky130_fd_sc_hd__o211a_1
X_15036_ _15483_/CLK _15036_/D _14073_/Y vssd1 vssd1 vccd1 vccd1 _15036_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12179_ _12240_/B _12179_/B vssd1 vssd1 vccd1 vccd1 _12181_/C sky130_fd_sc_hd__nand2_1
XFILLER_123_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater782_A _15615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08410_ _08388_/B _08410_/B vssd1 vssd1 vccd1 vccd1 _08639_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09390_ _09390_/A _09390_/B _09390_/C vssd1 vssd1 vccd1 vccd1 _09392_/A sky130_fd_sc_hd__and3_1
X_08341_ _08310_/A _08308_/A _08339_/X _08340_/X vssd1 vssd1 vccd1 vccd1 _08341_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ _08272_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14416__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__B _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput420 output420/A vssd1 vssd1 vccd1 vccd1 y_r_1[16] sky130_fd_sc_hd__buf_2
XFILLER_145_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput431 output431/A vssd1 vssd1 vccd1 vccd1 y_r_2[10] sky130_fd_sc_hd__buf_2
Xoutput442 output442/A vssd1 vssd1 vccd1 vccd1 y_r_2[5] sky130_fd_sc_hd__buf_2
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput453 output453/A vssd1 vssd1 vccd1 vccd1 y_r_3[15] sky130_fd_sc_hd__buf_2
Xoutput464 _15814_/X vssd1 vssd1 vccd1 vccd1 y_r_4[0] sky130_fd_sc_hd__buf_2
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput475 output475/A vssd1 vssd1 vccd1 vccd1 y_r_4[4] sky130_fd_sc_hd__buf_2
XFILLER_154_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput486 output486/A vssd1 vssd1 vccd1 vccd1 y_r_5[14] sky130_fd_sc_hd__buf_2
Xoutput497 _15619_/Q vssd1 vssd1 vccd1 vccd1 y_r_5[9] sky130_fd_sc_hd__buf_2
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14151__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_444 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07987_ _11435_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08005_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13990__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _09733_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _15309_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07522__A1 input100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _12630_/A _12803_/A vssd1 vssd1 vccd1 vccd1 _08732_/A sky130_fd_sc_hd__nor2_1
X_09588_ _15439_/Q _15423_/Q vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__or2b_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08728_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__nand2_1
XFILLER_179_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15132__D _15132_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _11550_/A _11550_/B vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__xor2_1
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _10501_/A _10501_/B vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__nand2_1
XFILLER_155_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14971__D _14971_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ _11687_/A _08157_/A _11480_/X vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14326__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input196_A x_r_4[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_689 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ _13220_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _14953_/D sky130_fd_sc_hd__xor2_2
XFILLER_183_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_970 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__A1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13151_ _13223_/B _13150_/C _13150_/A vssd1 vssd1 vccd1 vccd1 _13152_/B sky130_fd_sc_hd__o21ai_1
X_10363_ _10363_/A vssd1 vssd1 vccd1 vccd1 _15788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_833 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ _12102_/A vssd1 vssd1 vccd1 vccd1 _15586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _13192_/B _13082_/B vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input57_A x_i_3[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10437_/A _10294_/B vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _12308_/S _12231_/A _12228_/A vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__and3_1
XANTENNA__14061__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__A2 _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A1 _07761_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13984_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13984_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08994__A _15369_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15723_ _15725_/CLK _15723_/D _14799_/Y vssd1 vssd1 vccd1 vccd1 _15723_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A2 _15512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12935_ _12993_/A _12993_/B vssd1 vssd1 vccd1 vccd1 _12991_/B sky130_fd_sc_hd__xnor2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ _15689_/CLK _15654_/D _14727_/Y vssd1 vssd1 vccd1 vccd1 _15654_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ _12967_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__xnor2_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14605_/Y sky130_fd_sc_hd__inv_2
X_11817_ _11817_/A _11817_/B _11817_/C vssd1 vssd1 vccd1 vccd1 _11818_/B sky130_fd_sc_hd__nand3_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15585_ _15617_/CLK _15585_/D _14654_/Y vssd1 vssd1 vccd1 vccd1 _15585_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_973 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12797_ _12868_/B _12797_/B vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__xnor2_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15042__D _15042_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14536_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11749_/C sky130_fd_sc_hd__xnor2_1
XFILLER_109_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14467_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14467_/Y sky130_fd_sc_hd__inv_2
X_11679_ _11680_/A _11680_/B _11680_/C vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14236__A _14238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ _13416_/A _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__a21bo_1
XFILLER_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14398_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14398_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _13345_/A _13345_/B _13348_/X vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__a21o_2
XANTENNA__09049__B _15378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12325__A1 _12308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15439_/CLK _15019_/D _14055_/Y vssd1 vssd1 vccd1 vccd1 _15019_/Q sky130_fd_sc_hd__dfrtp_1
X_07910_ _15365_/Q _15349_/Q vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__nand2_1
X_08890_ _08890_/A _08959_/A vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__or2_1
XFILLER_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07841_ _07841_/A vssd1 vssd1 vccd1 vccd1 _15347_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater901 repeater902/X vssd1 vssd1 vccd1 vccd1 _07734_/A1 sky130_fd_sc_hd__buf_4
Xrepeater912 input200/X vssd1 vssd1 vccd1 vccd1 _07840_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater923 input186/X vssd1 vssd1 vccd1 vccd1 repeater923/X sky130_fd_sc_hd__buf_2
XFILLER_110_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater934 repeater935/X vssd1 vssd1 vccd1 vccd1 _07808_/A1 sky130_fd_sc_hd__buf_4
Xrepeater945 input153/X vssd1 vssd1 vccd1 vccd1 _07740_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07772_ _07772_/A vssd1 vssd1 vccd1 vccd1 _15381_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater956 input140/X vssd1 vssd1 vccd1 vccd1 _07894_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater967 repeater968/X vssd1 vssd1 vccd1 vccd1 _07408_/A1 sky130_fd_sc_hd__buf_4
XFILLER_204_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater978 repeater979/X vssd1 vssd1 vccd1 vccd1 _07524_/A1 sky130_fd_sc_hd__buf_4
X_09511_ _09511_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _15258_/D sky130_fd_sc_hd__xnor2_1
XFILLER_140_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07504__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09442_ _15533_/Q _15517_/Q vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09373_ _09371_/A _09371_/B _09372_/X vssd1 vssd1 vccd1 vccd1 _09375_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08324_ _08324_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08255_ _08289_/A _08288_/B _08255_/C vssd1 vssd1 vccd1 vccd1 _08307_/A sky130_fd_sc_hd__nor3_1
XFILLER_137_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14146__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _12144_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08190_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13985__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput261 output261/A vssd1 vssd1 vccd1 vccd1 y_i_0[10] sky130_fd_sc_hd__buf_2
Xoutput272 output272/A vssd1 vssd1 vccd1 vccd1 y_i_0[5] sky130_fd_sc_hd__buf_2
Xoutput283 _15658_/Q vssd1 vssd1 vccd1 vccd1 y_i_1[15] sky130_fd_sc_hd__buf_2
XFILLER_58_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput294 output294/A vssd1 vssd1 vccd1 vccd1 y_i_2[0] sky130_fd_sc_hd__buf_2
XFILLER_43_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_47 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ _15059_/Q _15092_/Q vssd1 vssd1 vccd1 vccd1 _09709_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10981_ _15173_/Q _15272_/Q vssd1 vssd1 vccd1 vccd1 _10982_/C sky130_fd_sc_hd__or2b_1
XANTENNA__08299__A2 _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input111_A x_i_6[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _12811_/A _12811_/B vssd1 vssd1 vccd1 vccd1 _12721_/B sky130_fd_sc_hd__xor2_1
XFILLER_74_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input209_A x_r_4[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__A _15726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ _08661_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__and2b_1
XFILLER_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ _11602_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nor2_1
X_12582_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _15679_/D sky130_fd_sc_hd__xnor2_1
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _15374_/CLK _15370_/D _14426_/Y vssd1 vssd1 vccd1 vccd1 _15370_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12783__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _14339_/A vssd1 vssd1 vccd1 vccd1 _14321_/Y sky130_fd_sc_hd__inv_2
X_11533_ _11531_/Y _11454_/B _11532_/X vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__o21a_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__A _14058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_947 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _11464_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__or2b_1
X_14252_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08054__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13203_ _13203_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _13203_/X sky130_fd_sc_hd__and2_1
X_10415_ _10415_/A vssd1 vssd1 vccd1 vccd1 _14947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14183_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14183_/Y sky130_fd_sc_hd__inv_2
X_11395_ _10194_/Y _11394_/B _10196_/B vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__o21ai_1
XFILLER_178_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08989__A _15368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10347_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _15786_/D sky130_fd_sc_hd__xor2_1
X_13134_ _15765_/Q _13558_/B vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__xor2_2
XFILLER_98_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _15764_/Q _13066_/B vssd1 vssd1 vccd1 vccd1 _13138_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10277_ _10277_/A vssd1 vssd1 vccd1 vccd1 _15771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08501__B _12688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _11940_/A _11940_/B _11951_/Y _11952_/Y _12454_/B vssd1 vssd1 vccd1 vccd1
+ _12223_/A sky130_fd_sc_hd__o311a_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output330_A output330/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07734__A1 _07734_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15037__D _15037_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output428_A _15585_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07832__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13967_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13967_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater578_A repeater579/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07498__A0 _15515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _15706_/CLK _15706_/D _14781_/Y vssd1 vssd1 vccd1 vccd1 _15706_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12918_ _12918_/A _13541_/A vssd1 vssd1 vccd1 vccd1 _15630_/D sky130_fd_sc_hd__xor2_4
XFILLER_59_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _13897_/A _13897_/C _13897_/B vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__o21a_1
XFILLER_179_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15637_ _15724_/CLK _15637_/D _14709_/Y vssd1 vssd1 vccd1 vccd1 _15637_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12849_ _12845_/A _13537_/A _12845_/B _12848_/Y vssd1 vssd1 vccd1 vccd1 _12918_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater745_A repeater746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _15568_/CLK _15568_/D _14635_/Y vssd1 vssd1 vccd1 vccd1 _15568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14519_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14519_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater912_A input200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15499_ _15528_/CLK _15499_/D _14563_/Y vssd1 vssd1 vccd1 vccd1 _15499_/Q sky130_fd_sc_hd__dfrtp_4
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A2 _11348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _09991_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _14931_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08942_ _08942_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _15188_/D sky130_fd_sc_hd__xnor2_1
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08873_ _15467_/Q _15451_/Q vssd1 vssd1 vccd1 vccd1 _08874_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater720 _15699_/Q vssd1 vssd1 vccd1 vccd1 output393/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07824_ _15355_/Q input175/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07825_/A sky130_fd_sc_hd__mux2_1
Xrepeater731 _15676_/Q vssd1 vssd1 vccd1 vccd1 output318/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater742 repeater743/X vssd1 vssd1 vccd1 vccd1 output282/A sky130_fd_sc_hd__buf_4
XFILLER_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater753 _15649_/Q vssd1 vssd1 vccd1 vccd1 output290/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater764 _15637_/Q vssd1 vssd1 vccd1 vccd1 output517/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07742__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater775 _15622_/Q vssd1 vssd1 vccd1 vccd1 output484/A sky130_fd_sc_hd__clkbuf_2
X_07755_ _15389_/Q _07755_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__mux2_1
Xrepeater786 _15606_/Q vssd1 vssd1 vccd1 vccd1 output450/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater797 _15594_/Q vssd1 vssd1 vccd1 vccd1 repeater797/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _07686_/A vssd1 vssd1 vccd1 vccd1 _15423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09425_ _09501_/A _09420_/B _09424_/X vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09035__B_N _15376_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09356_/A _09356_/B vssd1 vssd1 vccd1 vccd1 _15137_/D sky130_fd_sc_hd__nor2_1
XFILLER_139_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_740 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08307_ _08307_/A _08307_/B vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__or2_1
XFILLER_166_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _09285_/Y _09287_/B vssd1 vssd1 vccd1 vccd1 _09359_/A sky130_fd_sc_hd__nand2b_1
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _08243_/A _08225_/C _11842_/C vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__07661__A0 _15435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08169_ _08169_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14604__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ _15072_/Q _15237_/Q vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__or2_1
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _15025_/Q _15747_/Q vssd1 vssd1 vccd1 vccd1 _11181_/C sky130_fd_sc_hd__or2b_1
XFILLER_133_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08602__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10131_ _15142_/Q _15307_/Q vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09417__B _15512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input159_A x_r_1[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _15211_/Q _15112_/Q vssd1 vssd1 vccd1 vccd1 _10062_/X sky130_fd_sc_hd__and2_1
XFILLER_47_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07716__A1 _07716_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14870_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13821_ _13818_/A _13819_/A _13818_/B _13820_/Y vssd1 vssd1 vccd1 vccd1 _13822_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_85_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ _13752_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13753_/A sky130_fd_sc_hd__or2_1
X_10964_ _15152_/Q _10963_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10966_/C sky130_fd_sc_hd__a21o_1
XFILLER_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08049__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ _12703_/A _12703_/B _12703_/C vssd1 vssd1 vccd1 vccd1 _13022_/A sky130_fd_sc_hd__nand3_2
XFILLER_91_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13683_ _14975_/Q _13824_/B vssd1 vssd1 vccd1 vccd1 _13822_/A sky130_fd_sc_hd__xnor2_1
X_10895_ _10895_/A _11115_/A _10895_/C vssd1 vssd1 vccd1 vccd1 _10897_/A sky130_fd_sc_hd__and3_1
XFILLER_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15422_ _15699_/CLK _15422_/D _14482_/Y vssd1 vssd1 vccd1 vccd1 _15422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12634_ _12630_/A _08384_/C _08654_/A _12632_/Y _12813_/B vssd1 vssd1 vccd1 vccd1
+ _12635_/B sky130_fd_sc_hd__o221a_1
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15353_ _15477_/CLK _15353_/D _14408_/Y vssd1 vssd1 vccd1 vccd1 _15353_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13402__B _13576_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ _12268_/C _12563_/B _12564_/X vssd1 vssd1 vccd1 vccd1 _12566_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14304_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14304_/Y sky130_fd_sc_hd__inv_2
X_11516_ _11515_/Y _07995_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__mux2_1
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15284_ _15399_/CLK _15284_/D _14335_/Y vssd1 vssd1 vccd1 vccd1 _15284_/Q sky130_fd_sc_hd__dfrtp_4
X_12496_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output280_A output280/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output378_A _11121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14235_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14235_/Y sky130_fd_sc_hd__inv_2
X_11447_ _11658_/A _11447_/B _11447_/C vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__or3_1
XFILLER_153_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14514__A _14520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14166_/Y sky130_fd_sc_hd__inv_2
X_11378_ _15753_/Q _15031_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__a21o_1
XFILLER_153_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10329_ _10327_/Y _10329_/B vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__and2b_1
XFILLER_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13034_/A _13034_/B _13116_/X vssd1 vssd1 vccd1 vccd1 _13118_/B sky130_fd_sc_hd__a21oi_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12034__A _12178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14097_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14097_/Y sky130_fd_sc_hd__inv_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _12969_/B _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__and2b_1
XFILLER_117_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater695_A _14861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14999_ _15483_/CLK _14999_/D _14033_/Y vssd1 vssd1 vccd1 vccd1 _14999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_80_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07575_/S sky130_fd_sc_hd__buf_6
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07471_ _15528_/Q _07471_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_982 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _15576_/Q _15556_/Q vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__nor2_1
XFILLER_210_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_95_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09141_ _09136_/A _09140_/B _09136_/B vssd1 vssd1 vccd1 vccd1 _15234_/D sky130_fd_sc_hd__o21ba_1
XFILLER_194_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09072_/A _09072_/B vssd1 vssd1 vccd1 vccd1 _15219_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__xor2_1
XFILLER_194_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14424__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08422__A _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09872_/Y _09973_/B _09874_/B vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_33_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08925_/A _08925_/B _08973_/A vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__nor3_1
XFILLER_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08856_ _08855_/A _08855_/B _08939_/A vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__o21a_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _09253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater550 _11292_/X vssd1 vssd1 vccd1 vccd1 repeater550/X sky130_fd_sc_hd__buf_2
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater561 _11337_/X vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__clkbuf_2
X_07807_ _07807_/A vssd1 vssd1 vccd1 vccd1 _15364_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater572 _11079_/X vssd1 vssd1 vccd1 vccd1 repeater572/X sky130_fd_sc_hd__buf_2
Xrepeater583 _11197_/Y vssd1 vssd1 vccd1 vccd1 output513/A sky130_fd_sc_hd__clkbuf_2
X_08787_ _13885_/A _08782_/B _08786_/X vssd1 vssd1 vccd1 vccd1 _08788_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_48_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater594 _11367_/Y vssd1 vssd1 vccd1 vccd1 output445/A sky130_fd_sc_hd__buf_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _15397_/Q _07738_/A1 _07750_/S vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07669_ _15431_/Q _07669_/A1 _07697_/S vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09871__A1 _15185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09408_ _15510_/Q _15526_/Q vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__and2b_1
XFILLER_71_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10680_ _10999_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _15046_/D sky130_fd_sc_hd__xnor2_4
XFILLER_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09339_ _15411_/Q _15395_/Q vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__xor2_4
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07634__A0 _15448_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12573_/A sky130_fd_sc_hd__xnor2_2
XFILLER_126_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _10861_/Y _14987_/Q _11021_/B vssd1 vssd1 vccd1 vccd1 _11303_/C sky130_fd_sc_hd__a21o_1
XFILLER_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12281_ _12254_/A _12254_/B _12253_/A vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__a21o_1
XFILLER_107_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14334__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07647__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ _11230_/X _11235_/B vssd1 vssd1 vccd1 vccd1 _11232_/X sky130_fd_sc_hd__and2b_1
X_14020_ _14037_/A vssd1 vssd1 vccd1 vccd1 _14020_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11163_ _15746_/Q _15024_/Q vssd1 vssd1 vccd1 vccd1 _11163_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10814_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _15795_/D sky130_fd_sc_hd__xnor2_2
XFILLER_110_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _11093_/A _11093_/B _11348_/A vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12789__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _15184_/CLK _14922_/D _13952_/Y vssd1 vssd1 vccd1 vccd1 _14922_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ _10406_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _14977_/D sky130_fd_sc_hd__xnor2_1
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07382__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14853_/Y sky130_fd_sc_hd__inv_2
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13804_/A _13804_/B vssd1 vssd1 vccd1 vccd1 _13805_/B sky130_fd_sc_hd__xnor2_1
XFILLER_205_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14784_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11996_ _11994_/X _11996_/B vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__and2b_1
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13735_ _13723_/A _13725_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13740_/C sky130_fd_sc_hd__a21o_1
XFILLER_189_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _10945_/X _10950_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__and2b_2
XFILLER_16_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14509__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13666_ _13663_/A _13815_/A _13663_/B _13665_/X vssd1 vssd1 vccd1 vccd1 _13674_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10878_ _14958_/Q _14892_/Q vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output495_A _15617_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15405_ _15588_/CLK _15405_/D _14464_/Y vssd1 vssd1 vccd1 vccd1 _15405_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12615_/Y _12510_/B _12616_/Y vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__o21ai_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
X_13597_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _15089_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__15050__D _15050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_581 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15336_ _15725_/CLK _15336_/D _14390_/Y vssd1 vssd1 vccd1 vccd1 _15336_/Q sky130_fd_sc_hd__dfrtp_4
X_12548_ _12548_/A _12548_/B vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater610_A _11115_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15267_ _15268_/CLK _15267_/D _14317_/Y vssd1 vssd1 vccd1 vccd1 _15267_/Q sky130_fd_sc_hd__dfrtp_1
X_12479_ _12479_/A _12599_/A vssd1 vssd1 vccd1 vccd1 _12479_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14244__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater708_A _07536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07557__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14218_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15198_ _15472_/CLK _15198_/D _14245_/Y vssd1 vssd1 vccd1 vccd1 _15198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14149_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_791 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11807__S _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _08710_/X sky130_fd_sc_hd__or2_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ _15055_/Q _15088_/Q vssd1 vssd1 vccd1 vccd1 _09690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08641_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08641_/X sky130_fd_sc_hd__and2_1
XFILLER_6_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ _08728_/A _12970_/A vssd1 vssd1 vccd1 vccd1 _08615_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_1029 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12988__A1 _12910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__B2 _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _07523_/A vssd1 vssd1 vccd1 vccd1 _15503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14419__A _14419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07454_ _07454_/A vssd1 vssd1 vccd1 vccd1 _15537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08417__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ _07385_/A vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08136__B _08292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _15505_/Q _15489_/Q vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__xor2_2
XFILLER_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11778__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ _15379_/Q _15363_/Q vssd1 vssd1 vccd1 vccd1 _13628_/A sky130_fd_sc_hd__xnor2_1
XFILLER_191_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14154__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07467__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__xnor2_1
XFILLER_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13993__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07991__A _11458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_998 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09957_ _15199_/Q _15232_/Q vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__xor2_2
XFILLER_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08908_ _08907_/A _08907_/B _08963_/A vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _15221_/Q _15188_/Q vssd1 vssd1 vccd1 vccd1 _09889_/C sky130_fd_sc_hd__or2b_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _15348_/Q _15332_/Q vssd1 vssd1 vccd1 vccd1 _08841_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11849_/Y _11742_/A _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11852_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__B _12055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__nor2_2
XFILLER_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14974__D _14974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ _11824_/B _11781_/B vssd1 vssd1 vccd1 vccd1 _12403_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09844__A1 _15061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14329__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13520_ _13510_/A _13791_/B _13519_/Y vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__o21a_1
XFILLER_82_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10732_ _10728_/A _10725_/Y _10727_/B vssd1 vssd1 vccd1 vccd1 _10733_/B sky130_fd_sc_hd__o21ai_4
XFILLER_40_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10576__B _15298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ _13451_/A _15770_/Q vssd1 vssd1 vccd1 vccd1 _13480_/C sky130_fd_sc_hd__or2b_1
XFILLER_186_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ _10655_/Y _10659_/B _10657_/B vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__o21ai_4
XFILLER_16_1132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12402_ _12381_/B _12381_/C _12381_/D _12391_/B _12381_/A vssd1 vssd1 vccd1 vccd1
+ _12406_/B sky130_fd_sc_hd__a311o_1
XFILLER_185_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10594_ _10594_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _14990_/D sky130_fd_sc_hd__xnor2_1
X_13382_ _13438_/A _13381_/Y _13325_/A _13324_/A _13322_/B vssd1 vssd1 vccd1 vccd1
+ _13384_/B sky130_fd_sc_hd__o32a_1
XANTENNA_input87_A x_i_5[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _15279_/CLK _15121_/D _14163_/Y vssd1 vssd1 vccd1 vccd1 _15121_/Q sky130_fd_sc_hd__dfrtp_1
X_12333_ _12511_/A vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__inv_2
XANTENNA__09228__A_N _15496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14064__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_8
X_15052_ _15693_/CLK _15052_/D _14090_/Y vssd1 vssd1 vccd1 vccd1 _15052_/Q sky130_fd_sc_hd__dfrtp_4
X_12264_ _12214_/A _12218_/B _12214_/B vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21ba_1
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _14003_/A vssd1 vssd1 vccd1 vccd1 _14003_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ _11215_/A _11223_/A vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__nand2_1
X_12195_ _12132_/S _12204_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12195_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11146_ _11153_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11353_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11077_ _11077_/A _11077_/B _11344_/A vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__and3_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08335__A1 _11658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput150 x_r_1[12] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput161 x_r_1[8] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__clkbuf_1
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput172 x_r_2[3] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_hd__clkbuf_2
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08335__B2 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ _15399_/CLK _14905_/D _13934_/Y vssd1 vssd1 vccd1 vccd1 _14905_/Q sky130_fd_sc_hd__dfrtp_1
X_10028_ _10026_/Y _10028_/B vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__and2b_1
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput183 x_r_3[13] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__clkbuf_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output410_A output410/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output508_A output508/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput194 x_r_3[9] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15045__D _15045_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__B_N _15186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14836_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14836_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07840__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14767_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14767_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater560_A _11382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11979_ _11980_/A _11980_/B _11978_/Y vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__14239__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _13718_/A _13718_/B _13718_/C vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__nand3_1
XFILLER_189_475 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14698_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14698_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ _13649_/A _13649_/B vssd1 vssd1 vccd1 vccd1 _13651_/A sky130_fd_sc_hd__and2_1
XFILLER_158_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11598__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15319_ _15428_/CLK _15319_/D _14372_/Y vssd1 vssd1 vccd1 vccd1 _15319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_120_clk clkbuf_4_9_0_clk/X vssd1 vssd1 vccd1 vccd1 _15472_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09068__A _15478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09811_ _15443_/Q _15427_/Q _09810_/X vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10381__A1 _15086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _15098_/Q _15065_/Q vssd1 vssd1 vccd1 vccd1 _09743_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11764__C _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09673_ _15574_/Q _15554_/Q vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__or2b_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08624_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07750__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08555_ _08579_/B _08555_/B vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14149__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07506_ _15511_/Q input27/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08147__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08486_ _08486_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08548_/A sky130_fd_sc_hd__xor2_2
XFILLER_210_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13988__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ _15545_/Q _07437_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07438_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12892__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07986__A _15792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__A2 _12204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09107_ _15501_/Q _15485_/Q _09103_/B vssd1 vssd1 vccd1 vccd1 _09107_/X sky130_fd_sc_hd__o21a_1
XFILLER_202_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_111_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _15708_/CLK sky130_fd_sc_hd__clkbuf_16
X_09038_ _09038_/A _09038_/B _13618_/A vssd1 vssd1 vccd1 vccd1 _09038_/X sky130_fd_sc_hd__and3_1
XFILLER_191_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14612__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11000_ _10999_/B _10999_/C _10999_/A vssd1 vssd1 vccd1 vccd1 _11003_/C sky130_fd_sc_hd__a21o_1
XFILLER_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14969__D _14969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08610__A _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input141_A x_r_0[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input239_A x_r_6[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12951_ _12959_/A _12951_/B _12951_/C vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__or3_1
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11902_/A vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__inv_2
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ _15670_/CLK _15670_/D _14744_/Y vssd1 vssd1 vccd1 vccd1 _15670_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12882_/A _12882_/B vssd1 vssd1 vccd1 vccd1 _12902_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09119__B_N _15488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A vssd1 vssd1 vccd1 vccd1 _14640_/A sky130_fd_sc_hd__buf_12
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11833_ _11833_/A _11833_/B vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__or2_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__A _14219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14552_/Y sky130_fd_sc_hd__inv_2
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ _11764_/A _11797_/A _11876_/A vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__and3_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08057__A _08290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ _13494_/A _13782_/B _13502_/X vssd1 vssd1 vccd1 vccd1 _13510_/A sky130_fd_sc_hd__a21oi_2
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10713_/A _11014_/A _10714_/Y vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__o21ai_2
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14483_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09050__A_N _15378_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11695_ _11832_/A _11707_/A vssd1 vssd1 vccd1 vccd1 _11696_/B sky130_fd_sc_hd__nand2_1
XFILLER_186_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13377__A1 _13438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ _13431_/B _13433_/Y _13378_/B vssd1 vssd1 vccd1 vccd1 _13435_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10646_ _15271_/Q _15172_/Q vssd1 vssd1 vccd1 vccd1 _10647_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_871 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13365_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13425_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_831 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _15081_/CLK sky130_fd_sc_hd__clkbuf_16
X_10577_ _10577_/A _10577_/B _10622_/A vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__and3_1
XFILLER_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ _15367_/CLK _15104_/D _14145_/Y vssd1 vssd1 vccd1 vccd1 _15104_/Q sky130_fd_sc_hd__dfrtp_1
X_12316_ _12493_/A _12295_/B _12315_/X vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__a21oi_2
XFILLER_127_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13296_ _13290_/X _13723_/B _13291_/X _13294_/X _13295_/X vssd1 vssd1 vccd1 vccd1
+ _13345_/A sky130_fd_sc_hd__a311o_2
XANTENNA_output458_A output458/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15035_ _15509_/CLK _15035_/D _14072_/Y vssd1 vssd1 vccd1 vccd1 _15035_/Q sky130_fd_sc_hd__dfrtp_2
X_12247_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12247_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14522__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_902 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12178_ _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__or2_1
XFILLER_25_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08520__A _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11129_ _11129_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater775_A _15622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14819_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14819_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater942_A input159/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ _15799_/CLK _15799_/D _14879_/Y vssd1 vssd1 vccd1 vccd1 _15799_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08340_ _08310_/A _08308_/A _08328_/Y _08289_/X vssd1 vssd1 vccd1 vccd1 _08340_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08271_ _08271_/A _08271_/B vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_802 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput410 output410/A vssd1 vssd1 vccd1 vccd1 y_r_0[7] sky130_fd_sc_hd__buf_2
XFILLER_69_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput421 output421/A vssd1 vssd1 vccd1 vccd1 y_r_1[1] sky130_fd_sc_hd__buf_2
XFILLER_172_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput432 output432/A vssd1 vssd1 vccd1 vccd1 y_r_2[11] sky130_fd_sc_hd__buf_2
XFILLER_160_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput443 output443/A vssd1 vssd1 vccd1 vccd1 y_r_2[6] sky130_fd_sc_hd__buf_2
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14432__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput454 _15610_/Q vssd1 vssd1 vccd1 vccd1 y_r_3[16] sky130_fd_sc_hd__buf_2
Xoutput465 _11286_/X vssd1 vssd1 vccd1 vccd1 y_r_4[10] sky130_fd_sc_hd__buf_2
XANTENNA__08547__A1 _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput476 output476/A vssd1 vssd1 vccd1 vccd1 y_r_4[5] sky130_fd_sc_hd__buf_2
XFILLER_160_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput487 output487/A vssd1 vssd1 vccd1 vccd1 y_r_5[15] sky130_fd_sc_hd__buf_2
Xoutput498 _15816_/X vssd1 vssd1 vccd1 vccd1 y_r_6[0] sky130_fd_sc_hd__buf_2
XFILLER_113_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07986_ _15792_/Q vssd1 vssd1 vccd1 vccd1 _08290_/B sky130_fd_sc_hd__buf_12
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ _15062_/Q _15095_/Q vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__nand2_1
XFILLER_170_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12887__A _13366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09656_ _09656_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__and2_1
XFILLER_27_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09261__A _15505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _12881_/A vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__clkinv_2
XFILLER_103_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09587_ _15423_/Q _15439_/Q vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__or2b_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _12688_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08539_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08469_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__xor2_2
XANTENNA__14607__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _15254_/Q _15287_/Q vssd1 vssd1 vccd1 vccd1 _10501_/B sky130_fd_sc_hd__nand2_1
X_11480_ _11480_/A _11617_/A _11491_/A vssd1 vssd1 vccd1 vccd1 _11480_/X sky130_fd_sc_hd__and3_1
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10431_ _10430_/A _10430_/B _10086_/B vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__a21o_1
XFILLER_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input189_A x_r_3[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_982 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ _13150_/A _13223_/B _13150_/C vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__or3_1
X_10362_ _10360_/X _10368_/A vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__and2b_1
XFILLER_128_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12101_ _12099_/X _12156_/A vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__and2b_1
XFILLER_2_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_845 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10293_ _15120_/Q _15153_/Q vssd1 vssd1 vccd1 vccd1 _10294_/B sky130_fd_sc_hd__or2b_1
X_13081_ _13183_/A _12893_/C _13273_/A vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14342__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12032_ _12308_/S _12228_/A _12231_/A vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12885__A3 _12881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13983_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13983_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15722_ _15722_/CLK _15722_/D _14798_/Y vssd1 vssd1 vccd1 vccd1 _15722_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12934_ _12934_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _12993_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15653_ _15688_/CLK _15653_/D _14726_/Y vssd1 vssd1 vccd1 vccd1 _15653_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12794_/A _12793_/B _12793_/A vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__o21bai_1
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13598__A1 _15368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14604_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14604_/Y sky130_fd_sc_hd__inv_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__A _15752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ _11817_/A _11817_/B _11817_/C vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__a21o_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15732_/CLK _15584_/D _14653_/Y vssd1 vssd1 vccd1 vccd1 _15584_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12796_ _12749_/A _12749_/B _12795_/Y vssd1 vssd1 vccd1 vccd1 _12797_/B sky130_fd_sc_hd__a21oi_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14538_/A vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__inv_2
X_11747_ _11906_/A _11696_/B _11701_/B _11746_/Y vssd1 vssd1 vccd1 vccd1 _11834_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14517__A _14517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13421__A _13422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14466_/Y sky130_fd_sc_hd__inv_2
X_11678_ _11678_/A _11678_/B vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__xnor2_1
XFILLER_144_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08515__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13417_ _13417_/A _13417_/B vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__or2_1
X_10629_ _15169_/Q _15268_/Q vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__or2b_1
XFILLER_139_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12037__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14397_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14397_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13348_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11876__A _11876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14252__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13279_ _13277_/X _13316_/B vssd1 vssd1 vccd1 vccd1 _13280_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07565__S _07579_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ _15439_/CLK _15018_/D _14054_/Y vssd1 vssd1 vccd1 vccd1 _15018_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_1191 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater892_A input231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1044 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07840_ _15347_/Q _07840_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07841_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09065__B _15364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater902 input219/X vssd1 vssd1 vccd1 vccd1 repeater902/X sky130_fd_sc_hd__buf_2
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater913 input20/X vssd1 vssd1 vccd1 vccd1 _07490_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_111_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater924 input185/X vssd1 vssd1 vccd1 vccd1 _07675_/A1 sky130_fd_sc_hd__buf_4
Xrepeater935 input168/X vssd1 vssd1 vccd1 vccd1 repeater935/X sky130_fd_sc_hd__buf_2
Xrepeater946 input152/X vssd1 vssd1 vccd1 vccd1 _07742_/A1 sky130_fd_sc_hd__buf_4
X_07771_ _15381_/Q _07771_/A1 _07795_/S vssd1 vssd1 vccd1 vccd1 _07772_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater957 input139/X vssd1 vssd1 vccd1 vccd1 _07896_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater968 input123/X vssd1 vssd1 vccd1 vccd1 repeater968/X sky130_fd_sc_hd__buf_2
XANTENNA__13825__A2 _13822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _09431_/Y _09509_/B _09433_/B vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__o21ai_1
Xrepeater979 input114/X vssd1 vssd1 vccd1 vccd1 repeater979/X sky130_fd_sc_hd__buf_2
XFILLER_65_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09441_ _15533_/Q _15517_/Q vssd1 vssd1 vccd1 vccd1 _09441_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15811__A _15811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ _15404_/Q _15388_/Q vssd1 vssd1 vccd1 vccd1 _09372_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08323_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__xor2_1
XFILLER_71_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14427__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ _08254_/A _08254_/B vssd1 vssd1 vccd1 vccd1 _08255_/C sky130_fd_sc_hd__xor2_1
XFILLER_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _08185_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14162__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput262 output262/A vssd1 vssd1 vccd1 vccd1 y_i_0[11] sky130_fd_sc_hd__buf_2
XANTENNA__07475__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput273 output273/A vssd1 vssd1 vccd1 vccd1 y_i_0[6] sky130_fd_sc_hd__buf_2
Xoutput284 output284/A vssd1 vssd1 vccd1 vccd1 y_i_1[16] sky130_fd_sc_hd__buf_2
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput295 _10927_/X vssd1 vssd1 vccd1 vccd1 y_i_2[10] sky130_fd_sc_hd__buf_2
XFILLER_134_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08940__A1 _15463_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _07969_/A _11248_/A vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09708_ _09830_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _15714_/D sky130_fd_sc_hd__xnor2_1
X_10980_ _10980_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10982_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13292__A3 _13713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ _09639_/A _09639_/B vssd1 vssd1 vccd1 vccd1 _15304_/D sky130_fd_sc_hd__xor2_1
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _08660_/B _12650_/B vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__and2b_1
XANTENNA_input104_A x_i_6[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11601_ _12228_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11602_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_911 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12581_ _12579_/Y _12578_/B _12580_/Y vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__o21ai_1
XFILLER_168_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14337__A _14339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14320_ _14420_/A vssd1 vssd1 vccd1 vccd1 _14339_/A sky130_fd_sc_hd__buf_8
XANTENNA__12783__C _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _11532_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__or2_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_999 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14251_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14251_/Y sky130_fd_sc_hd__inv_2
X_11463_ _11463_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _12360_/B sky130_fd_sc_hd__xnor2_4
XFILLER_183_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13274_/B _13202_/B vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__nand2_2
XFILLER_7_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10414_ _10414_/A _10417_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__and2_1
X_14182_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ _11394_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _15728_/D sky130_fd_sc_hd__xnor2_1
XFILLER_174_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11696__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ _13703_/B _13133_/B vssd1 vssd1 vccd1 vccd1 _13558_/B sky130_fd_sc_hd__xor2_4
XFILLER_180_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _15130_/Q _15163_/Q vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__xor2_2
XFILLER_139_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14072__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13504__A1 _13352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13290_/A _13700_/A vssd1 vssd1 vccd1 vccd1 _13066_/B sky130_fd_sc_hd__xnor2_1
X_10276_ _10274_/X _10279_/B vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12304__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _12439_/B _12427_/B vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__xor2_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14800__A _14801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output323_A output323/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13966_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13966_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1102 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10759__B _15784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07498__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15705_ _15705_/CLK _15705_/D _14780_/Y vssd1 vssd1 vccd1 vccd1 _15705_/Q sky130_fd_sc_hd__dfrtp_4
X_12917_ _13545_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__xnor2_4
XFILLER_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13897_ _13897_/A _13897_/B _13897_/C vssd1 vssd1 vccd1 vccd1 _13899_/A sky130_fd_sc_hd__nor3_1
XFILLER_98_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12848_ _12848_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nor2_1
X_15636_ _15768_/CLK _15636_/D _14708_/Y vssd1 vssd1 vccd1 vccd1 _15636_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15567_ _15569_/CLK _15567_/D _14634_/Y vssd1 vssd1 vccd1 vccd1 _15567_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_187_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12779_/A _12779_/B vssd1 vssd1 vccd1 vccd1 _12805_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_242 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14247__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14518_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14518_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15498_ _15498_/CLK _15498_/D _14562_/Y vssd1 vssd1 vccd1 vccd1 _15498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_908 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14449_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14449_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater905_A input214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1106 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07422__A1 _07422_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09990_ _09990_/A _09990_/B _09990_/C vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__and3_1
XFILLER_171_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ _15463_/Q _15447_/Q _08940_/X vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__a21o_1
XFILLER_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08872_ _15467_/Q _15451_/Q vssd1 vssd1 vccd1 vccd1 _08872_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14710__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater710 _07900_/S vssd1 vssd1 vccd1 vccd1 _07892_/S sky130_fd_sc_hd__buf_6
XANTENNA__09804__A _15441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater721 _15697_/Q vssd1 vssd1 vccd1 vccd1 output391/A sky130_fd_sc_hd__clkbuf_2
X_07823_ _07823_/A vssd1 vssd1 vccd1 vccd1 _15356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater732 repeater733/X vssd1 vssd1 vccd1 vccd1 output317/A sky130_fd_sc_hd__buf_6
XFILLER_111_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater743 _15657_/Q vssd1 vssd1 vccd1 vccd1 repeater743/X sky130_fd_sc_hd__buf_2
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater754 _15647_/Q vssd1 vssd1 vccd1 vccd1 output288/A sky130_fd_sc_hd__clkbuf_2
Xrepeater765 _15634_/Q vssd1 vssd1 vccd1 vccd1 output530/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13326__A _14920_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _07754_/A vssd1 vssd1 vccd1 vccd1 _15390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater776 repeater777/X vssd1 vssd1 vccd1 vccd1 output482/A sky130_fd_sc_hd__buf_4
XANTENNA__12230__A _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater787 repeater788/X vssd1 vssd1 vccd1 vccd1 output448/A sky130_fd_sc_hd__buf_4
Xrepeater798 _15593_/Q vssd1 vssd1 vccd1 vccd1 output420/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07685_ _15423_/Q input180/X _07687_/S vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_91_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _15346_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09424_ _15528_/Q _15512_/Q vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ _09354_/A _09354_/C _09354_/B vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14157__A _14158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ _08289_/A _08288_/B _08255_/C vssd1 vssd1 vccd1 vccd1 _08307_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _15400_/Q _15384_/Q vssd1 vssd1 vccd1 vccd1 _09287_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08237_ _08237_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07661__A1 input255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13996__A _13997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07994__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ _11928_/A _11832_/A vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__xor2_2
XFILLER_134_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08099_ _08328_/A _08286_/A vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__or2_1
XFILLER_69_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ _15142_/Q _15307_/Q vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__or2_1
XFILLER_134_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08829__A_N _15330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ _10417_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _14980_/D sky130_fd_sc_hd__xnor2_2
XFILLER_173_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14620__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14977__D _14977_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13820_ _14974_/Q _13820_/B vssd1 vssd1 vccd1 vccd1 _13820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input221_A x_r_5[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _14981_/Q _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13752_/B sky130_fd_sc_hd__and3b_1
XFILLER_84_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ _10963_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_82_clk _14904_/CLK vssd1 vssd1 vccd1 vccd1 _15782_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ _15760_/Q vssd1 vssd1 vccd1 vccd1 _12843_/A sky130_fd_sc_hd__inv_2
X_13682_ _13682_/A _13682_/B vssd1 vssd1 vccd1 vccd1 _13824_/B sky130_fd_sc_hd__xnor2_4
XFILLER_204_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ _14893_/Q _14959_/Q vssd1 vssd1 vccd1 vccd1 _10895_/C sky130_fd_sc_hd__or2b_1
XFILLER_43_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _15434_/CLK _15421_/D _14480_/Y vssd1 vssd1 vccd1 vccd1 _15421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_203_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12633_ _12881_/A _12921_/A vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__or2b_1
XFILLER_197_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14067__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ _15352_/CLK _15352_/D _14407_/Y vssd1 vssd1 vccd1 vccd1 _15352_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_184_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _15738_/Q _12564_/B vssd1 vssd1 vccd1 vccd1 _12564_/X sky130_fd_sc_hd__and2_1
XFILLER_129_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1076 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14303_/Y sky130_fd_sc_hd__inv_2
X_11515_ _11797_/A vssd1 vssd1 vccd1 vccd1 _11515_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15283_ _15399_/CLK _15283_/D _14334_/Y vssd1 vssd1 vccd1 vccd1 _15283_/Q sky130_fd_sc_hd__dfrtp_4
X_12495_ _14951_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_767 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14234_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14234_/Y sky130_fd_sc_hd__inv_2
X_11446_ _11678_/A _11770_/A vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_610 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output273_A output273/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__A1 _07404_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14165_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11377_ _11377_/A _11377_/B vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__nor2_2
X_13116_ _13033_/B _13116_/B vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__and2b_1
X_10328_ _15127_/Q _15160_/Q vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__nand2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14096_/Y sky130_fd_sc_hd__inv_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output440_A output440/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13124_/B _13047_/B vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__nand2_1
XFILLER_152_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10259_ _10259_/A _10267_/A vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14530__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater590_A _10912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater688_A _14269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14998_ _15498_/CLK _14998_/D _14032_/Y vssd1 vssd1 vccd1 vccd1 _14998_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_207_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13949_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13949_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07470_ _07470_/A vssd1 vssd1 vccd1 vccd1 _15529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15619_ _15689_/CLK _15619_/D _14690_/Y vssd1 vssd1 vccd1 vccd1 _15619_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ _09271_/A _09140_/B vssd1 vssd1 vccd1 vccd1 _15233_/D sky130_fd_sc_hd__xor2_1
XFILLER_147_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _15493_/Q _15477_/Q _09219_/C vssd1 vssd1 vccd1 vccd1 _09072_/B sky130_fd_sc_hd__and3_1
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14705__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08022_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _08023_/B sky130_fd_sc_hd__xor2_1
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_598 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08703__A _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08422__B _12810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _14923_/D sky130_fd_sc_hd__xnor2_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09148__A1 _15562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ _15475_/Q _15459_/Q vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14440__A _14842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07753__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _08855_/A _08855_/B _08939_/A vssd1 vssd1 vccd1 vccd1 _08857_/A sky130_fd_sc_hd__nor3_1
XFILLER_170_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater540 _10962_/Y vssd1 vssd1 vccd1 vccd1 output301/A sky130_fd_sc_hd__clkbuf_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater551 _11140_/Y vssd1 vssd1 vccd1 vccd1 output368/A sky130_fd_sc_hd__clkbuf_2
X_07806_ _15364_/Q input169/X _07856_/S vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__mux2_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater562 _11285_/X vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__clkbuf_2
X_08786_ _15338_/Q _15322_/Q vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__and2b_1
Xrepeater573 _10781_/X vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__buf_2
Xrepeater584 _11125_/Y vssd1 vssd1 vccd1 vccd1 output363/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater595 _11321_/Y vssd1 vssd1 vccd1 vccd1 output341/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _07737_/A vssd1 vssd1 vccd1 vccd1 _15398_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _15680_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07668_ _07668_/A vssd1 vssd1 vccd1 vccd1 _15432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ _15526_/Q _15510_/Q vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__and2b_1
XFILLER_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07882__A1 input146/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07599_ _07599_/A vssd1 vssd1 vccd1 vccd1 _15466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ _09336_/A _09397_/A _09337_/Y vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__o21ai_4
XFILLER_166_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07634__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _15507_/Q vssd1 vssd1 vccd1 vccd1 _09269_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14615__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _11300_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11300_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_154_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _12280_/A _12280_/B vssd1 vssd1 vccd1 vccd1 _12291_/A sky130_fd_sc_hd__xnor2_2
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _11230_/A _11230_/B _11382_/A vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__a21o_1
XANTENNA_input171_A x_r_2[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12135__A _12244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ _11357_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11167_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09139__A1 _15507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10113_ _10109_/A _10106_/Y _10108_/B vssd1 vssd1 vccd1 vccd1 _10114_/B sky130_fd_sc_hd__o21ai_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ _11093_/A _11093_/B _11348_/A vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__and3_1
XANTENNA__14350__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07663__S _07695_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12789__B _13220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A x_i_1[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ _15184_/CLK _14921_/D _13951_/Y vssd1 vssd1 vccd1 vccd1 _14921_/Q sky130_fd_sc_hd__dfrtp_2
X_10044_ _10036_/Y _10040_/B _10038_/B vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__o21ai_1
XFILLER_49_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13891__B1 _13890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14852_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ _13803_/A _13519_/B vssd1 vssd1 vccd1 vccd1 _13804_/A sky130_fd_sc_hd__or2b_1
XFILLER_21_1053 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14783_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14783_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ _12312_/S _12204_/A _11994_/B _11994_/C vssd1 vssd1 vccd1 vccd1 _11996_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15777_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _13718_/B _13718_/C _13725_/C _13718_/A vssd1 vssd1 vccd1 vccd1 _13740_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10946_ _10945_/A _10945_/B _11134_/A vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _14973_/Q _13816_/B vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__and2_1
XFILLER_143_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877_ _14958_/Q _14892_/Q vssd1 vssd1 vccd1 vccd1 _10877_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11214__A _15031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15411_/CLK _15404_/D _14463_/Y vssd1 vssd1 vccd1 vccd1 _15404_/Q sky130_fd_sc_hd__dfrtp_1
X_12616_ _12613_/A _12613_/B _12614_/A vssd1 vssd1 vccd1 vccd1 _12616_/Y sky130_fd_sc_hd__o21ai_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output390_A _15696_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13596_ _15367_/Q _15351_/Q _13595_/X vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__a21o_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output488_A output488/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15335_ _15428_/CLK _15335_/D _14389_/Y vssd1 vssd1 vccd1 vccd1 _15335_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_531 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12547_ _12547_/A _12548_/B vssd1 vssd1 vccd1 vccd1 _15617_/D sky130_fd_sc_hd__xor2_1
XFILLER_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14525__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15266_ _15268_/CLK _15266_/D _14316_/Y vssd1 vssd1 vccd1 vccd1 _15266_/Q sky130_fd_sc_hd__dfrtp_1
X_12478_ _12478_/A _12599_/A _12478_/C vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__nand3_1
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10772__B _15786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14217_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ _10287_/B _11427_/B _11428_/Y vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_repeater603_A _11051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15197_ _15472_/CLK _15197_/D _14244_/Y vssd1 vssd1 vccd1 vccd1 _15197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14148_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11884__A _12122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__buf_12
XANTENNA__14260__A _14420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07573__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater972_A repeater973/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08640_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08640_/X sky130_fd_sc_hd__or2_1
XFILLER_187_1013 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07561__A0 _15484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _13046_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _15435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _15503_/Q input100/X _07538_/S vssd1 vssd1 vccd1 vccd1 _07523_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07864__A1 _07864_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13323__B _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ _15537_/Q _07453_/A1 _07485_/S vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_819 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15241__D _15241_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__B _12921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_649 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07384_ _15575_/Q input120/X _07432_/S vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09123_ _09121_/A _09254_/B _09122_/X vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__a21o_1
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07616__A1 _07616_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10963__A _10963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14435__A _14435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__S _07750_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _09054_/A _09056_/B vssd1 vssd1 vccd1 vccd1 _15115_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10777__A_N _15787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08433__A _08728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08005_ _11458_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__nor2_1
XFILLER_194_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_602 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11794__A _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _09956_/A vssd1 vssd1 vccd1 vccd1 _14967_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14170__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07483__S _07485_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08907_ _08907_/A _08907_/B _08963_/A vssd1 vssd1 vccd1 vccd1 _08907_/X sky130_fd_sc_hd__and3_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09887_ _09885_/Y _09887_/B vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__and2b_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _15083_/D sky130_fd_sc_hd__nor2_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _15336_/Q _15320_/Q vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__xnor2_2
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _15803_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _15790_/Q _15724_/Q vssd1 vssd1 vccd1 vccd1 _10801_/B sky130_fd_sc_hd__and2b_1
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11685_/A _11685_/B _11681_/A vssd1 vssd1 vccd1 vccd1 _11781_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11960__C _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08608__A _12630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _10731_/A _10731_/B vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__nand2_2
XFILLER_14_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_638 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ _13452_/A _13579_/A vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__xor2_1
X_10662_ _10662_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__nand2_2
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _14943_/Q _12401_/B _12401_/C vssd1 vssd1 vccd1 vccd1 _12410_/C sky130_fd_sc_hd__and3_1
XFILLER_107_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13381_ _13390_/A _13381_/B vssd1 vssd1 vccd1 vccd1 _13381_/Y sky130_fd_sc_hd__nand2_1
X_10593_ _10493_/Y _10592_/B _10495_/B vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__14345__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _15792_/CLK _15120_/D _14162_/Y vssd1 vssd1 vccd1 vccd1 _15120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12332_ _12332_/A _12332_/B vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__xnor2_4
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15051_ _15693_/CLK _15051_/D _14089_/Y vssd1 vssd1 vccd1 vccd1 _15051_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _12261_/X _12263_/B vssd1 vssd1 vccd1 vccd1 _12484_/A sky130_fd_sc_hd__and2b_1
XFILLER_126_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _14003_/A vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__inv_2
X_11214_ _15031_/Q _15753_/Q vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__or2b_1
X_12194_ _12252_/A _12194_/B vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__or2_1
XFILLER_123_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11145_ _15743_/Q _15021_/Q vssd1 vssd1 vccd1 vccd1 _11146_/B sky130_fd_sc_hd__or2b_1
XANTENNA__14080__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__A0 _15371_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_94_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__nor2_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 x_r_0[3] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_1
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput151 x_r_1[13] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_1
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14904_ _14904_/CLK _14904_/D _13933_/Y vssd1 vssd1 vccd1 vccd1 _14904_/Q sky130_fd_sc_hd__dfrtp_1
X_10027_ _15205_/Q _15106_/Q vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput162 x_r_1[9] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__buf_4
Xinput173 x_r_2[4] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07543__A0 _15493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput184 x_r_3[14] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput195 x_r_4[0] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_2
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14835_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output403_A output403/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15592_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _12056_/B _11978_/B vssd1 vssd1 vccd1 vccd1 _11978_/Y sky130_fd_sc_hd__nand2_1
X_14766_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14766_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ _14899_/Q _14965_/Q vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__or2b_1
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13717_ _13718_/B _13718_/C _13718_/A vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07846__A1 input197/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14697_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14697_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater553_A _11385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_32_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ _13648_/A _13648_/B vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__nand2_2
XFILLER_72_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11879__A _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater720_A _15699_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13579_ _13579_/A _13579_/B vssd1 vssd1 vccd1 vccd1 _15606_/D sky130_fd_sc_hd__xor2_1
XFILLER_185_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater818_A input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14255__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11598__B _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09349__A _15381_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ _15722_/CLK _15318_/D _14371_/Y vssd1 vssd1 vccd1 vccd1 _15318_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_47_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ _15249_/CLK _15249_/D _14298_/Y vssd1 vssd1 vccd1 vccd1 _15249_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09810_ _15443_/Q _15427_/Q _09809_/B vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10381__A2 _10380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _15065_/Q _15098_/Q vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__and2b_1
XFILLER_100_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_105_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15814__A _15814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _15313_/D sky130_fd_sc_hd__xor2_1
XANTENNA__07534__A0 _15497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_939 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_894 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ _08725_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _15444_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_950 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08550_/A _08550_/B _08553_/X vssd1 vssd1 vccd1 vccd1 _08555_/B sky130_fd_sc_hd__a21oi_1
XFILLER_78_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07505_ _07505_/A vssd1 vssd1 vccd1 vccd1 _15512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08485_ _13381_/B _08491_/B vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__xnor2_2
XFILLER_210_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08147__B _11687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07436_ _07436_/A vssd1 vssd1 vccd1 vccd1 _15546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10693__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14165__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _09113_/A _09114_/A vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__or2_1
XFILLER_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09037_ _09037_/A _09045_/A vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__nand2_1
XFILLER_201_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08610__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _09939_/A _09939_/B _09993_/A vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__and3_1
XFILLER_86_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_19_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _12871_/A _12871_/B _12949_/X vssd1 vssd1 vccd1 vccd1 _13054_/A sky130_fd_sc_hd__a21boi_4
XFILLER_46_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input134_A x_r_0[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11901_ _11901_/A _11901_/B _11901_/C vssd1 vssd1 vccd1 vccd1 _11902_/A sky130_fd_sc_hd__and3_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12881_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _12906_/B sky130_fd_sc_hd__nand2_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11832_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__nand2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14620_/Y sky130_fd_sc_hd__inv_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07828__A1 _07828_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14551_/Y sky130_fd_sc_hd__inv_2
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__inv_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__A1 _13201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _15282_/Q _15183_/Q vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nand2_1
X_13502_ _13790_/B _13790_/A vssd1 vssd1 vccd1 vccd1 _13502_/X sky130_fd_sc_hd__and2b_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14482_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11742_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11702_/A sky130_fd_sc_hd__nor2_1
XFILLER_186_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13433_ _13433_/A vssd1 vssd1 vccd1 vccd1 _13433_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13377__A2 _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ _15271_/Q _15172_/Q vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14075__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07388__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _13362_/X _13425_/A vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08073__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_883 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10576_ _15265_/Q _15298_/Q vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__xor2_2
XFILLER_6_843 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ _12291_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12315_/X sky130_fd_sc_hd__and2b_1
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _15367_/CLK _15103_/D _14144_/Y vssd1 vssd1 vccd1 vccd1 _15103_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295_ _13737_/B _13295_/B vssd1 vssd1 vccd1 vccd1 _13295_/X sky130_fd_sc_hd__and2_1
XANTENNA__14803__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15509_/CLK _15034_/D _14071_/Y vssd1 vssd1 vccd1 vccd1 _15034_/Q sky130_fd_sc_hd__dfrtp_4
X_12246_ _12247_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__and2_1
XFILLER_135_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_914 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08520__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11128_ _11127_/B _11127_/C _11127_/A vssd1 vssd1 vccd1 vccd1 _11129_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08012__S _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_958 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output520_A output520/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11059_ _11066_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__nand2_2
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater670_A _14709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater768_A _15630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13154__A _13390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14818_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14818_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15798_ _15799_/CLK _15798_/D _14878_/Y vssd1 vssd1 vccd1 vccd1 _15798_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ _14750_/A vssd1 vssd1 vccd1 vccd1 _14749_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08270_ _11499_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__xnor2_2
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09079__A _15496_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput400 _10790_/X vssd1 vssd1 vccd1 vccd1 y_r_0[13] sky130_fd_sc_hd__buf_2
XANTENNA__14713__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _15568_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput411 output411/A vssd1 vssd1 vccd1 vccd1 y_r_0[8] sky130_fd_sc_hd__buf_2
Xoutput422 _15579_/Q vssd1 vssd1 vccd1 vccd1 y_r_1[2] sky130_fd_sc_hd__buf_2
XFILLER_160_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput433 output433/A vssd1 vssd1 vccd1 vccd1 y_r_2[12] sky130_fd_sc_hd__buf_2
XFILLER_172_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput444 output444/A vssd1 vssd1 vccd1 vccd1 y_r_2[7] sky130_fd_sc_hd__buf_2
Xoutput455 output455/A vssd1 vssd1 vccd1 vccd1 y_r_3[1] sky130_fd_sc_hd__buf_2
XANTENNA__11548__S _11707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput466 output466/A vssd1 vssd1 vccd1 vccd1 y_r_4[11] sky130_fd_sc_hd__buf_2
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput477 _11269_/Y vssd1 vssd1 vccd1 vccd1 y_r_4[6] sky130_fd_sc_hd__buf_2
XFILLER_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput488 output488/A vssd1 vssd1 vccd1 vccd1 y_r_5[16] sky130_fd_sc_hd__buf_2
Xoutput499 _11212_/X vssd1 vssd1 vccd1 vccd1 y_r_6[10] sky130_fd_sc_hd__buf_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07985_ _11458_/A _08074_/C vssd1 vssd1 vccd1 vccd1 _08087_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09724_ _15062_/Q _15095_/Q vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__or2_1
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07761__S _07765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__B _13273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _09654_/B _09654_/C _09654_/A vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__o21ai_1
XFILLER_132_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08606_ _12810_/A _08603_/B _08500_/Y _12654_/A _08605_/X vssd1 vssd1 vccd1 vccd1
+ _08606_/X sky130_fd_sc_hd__a221o_1
X_09586_ _15438_/Q _15422_/Q vssd1 vssd1 vccd1 vccd1 _09590_/B sky130_fd_sc_hd__or2b_1
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_8
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08158__A _11832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13999__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08546_/A _08546_/B vssd1 vssd1 vccd1 vccd1 _08540_/A sky130_fd_sc_hd__xor2_2
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_975 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08468_ _08669_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__xnor2_2
XFILLER_204_1119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_755 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07419_/A vssd1 vssd1 vccd1 vccd1 _15554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _08441_/A _08399_/B _13201_/A vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__or3b_1
XFILLER_17_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12408__A _14944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10430_ _10430_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _14952_/D sky130_fd_sc_hd__xor2_2
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _10360_/A _10360_/B _10480_/A vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__a21o_1
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_994 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14623__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ _12099_/A _12099_/B _12553_/A vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__a21o_1
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13080_ _13357_/B vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__inv_2
X_10292_ _15153_/Q _15120_/Q vssd1 vssd1 vccd1 vccd1 _10437_/A sky130_fd_sc_hd__or2b_1
XFILLER_2_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_857 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ _12031_/A _12031_/B vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__or2_1
XFILLER_88_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input251_A x_r_7[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12143__A _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _13997_/A vssd1 vssd1 vccd1 vccd1 _13982_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07671__S _07697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15721_ _15722_/CLK _15721_/D _14797_/Y vssd1 vssd1 vccd1 vccd1 _15721_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _13203_/A _12933_/B _13006_/A _12931_/X vssd1 vssd1 vccd1 vccd1 _13006_/B
+ sky130_fd_sc_hd__or4bb_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15652_ _15687_/CLK _15652_/D _14725_/Y vssd1 vssd1 vccd1 vccd1 _15652_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ _12864_/A _12951_/C vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__xnor2_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14603_/Y sky130_fd_sc_hd__inv_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _11815_/A _11815_/B vssd1 vssd1 vccd1 vccd1 _11817_/C sky130_fd_sc_hd__nand2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_700 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15583_ _15617_/CLK _15583_/D _14652_/Y vssd1 vssd1 vccd1 vccd1 _15583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12795_ _12795_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12795_/Y sky130_fd_sc_hd__nor2_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11746_/Y sky130_fd_sc_hd__nand2_1
X_14534_ _14540_/A vssd1 vssd1 vccd1 vccd1 _14534_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_934 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11678_/B sky130_fd_sc_hd__xor2_1
X_14465_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14465_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__B _12871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13416_ _13416_/A _15052_/Q vssd1 vssd1 vccd1 vccd1 _13417_/B sky130_fd_sc_hd__nor2_1
X_10628_ _10628_/A _10628_/B vssd1 vssd1 vccd1 vccd1 _15003_/D sky130_fd_sc_hd__xnor2_1
XANTENNA_output470_A output470/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14396_ _14399_/A vssd1 vssd1 vccd1 vccd1 _14396_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_651 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13347_ _13347_/A _13403_/A vssd1 vssd1 vccd1 vccd1 _15636_/D sky130_fd_sc_hd__xnor2_1
XFILLER_183_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ _10558_/A _10558_/B _10612_/A vssd1 vssd1 vccd1 vccd1 _10565_/B sky130_fd_sc_hd__a21o_1
XFILLER_143_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14533__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07846__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A_N _15468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _13100_/A _13100_/B _13098_/A _13206_/Y _13208_/A vssd1 vssd1 vccd1 vccd1
+ _13316_/B sky130_fd_sc_hd__a311o_1
XANTENNA__08531__A _13319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15017_ _15435_/CLK _15017_/D _14053_/Y vssd1 vssd1 vccd1 vccd1 _15017_/Q sky130_fd_sc_hd__dfrtp_1
X_12229_ _12231_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13149__A _13491_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater903 input217/X vssd1 vssd1 vccd1 vccd1 _07708_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater885_A input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_243 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater914 input199/X vssd1 vssd1 vccd1 vccd1 _07842_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater925 input184/X vssd1 vssd1 vccd1 vccd1 _07677_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater936 input165/X vssd1 vssd1 vccd1 vccd1 _07814_/A1 sky130_fd_sc_hd__clkbuf_2
X_07770_ _07770_/A vssd1 vssd1 vccd1 vccd1 _15382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater947 input151/X vssd1 vssd1 vccd1 vccd1 _07744_/A1 sky130_fd_sc_hd__clkbuf_2
Xrepeater958 input137/X vssd1 vssd1 vccd1 vccd1 _07870_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07581__S _07591_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater969 input122/X vssd1 vssd1 vccd1 vccd1 _07410_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ _09511_/A _09440_/B vssd1 vssd1 vccd1 vccd1 _15274_/D sky130_fd_sc_hd__xor2_2
XFILLER_80_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _15142_/D sky130_fd_sc_hd__xor2_1
XFILLER_197_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14708__A _14714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__nand2_1
XFILLER_177_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08254_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12228__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _11687_/A _11491_/A vssd1 vssd1 vccd1 vccd1 _08185_/A sky130_fd_sc_hd__nand2_1
XFILLER_192_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14443__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_655 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput263 _11080_/X vssd1 vssd1 vccd1 vccd1 y_i_0[12] sky130_fd_sc_hd__buf_2
XFILLER_121_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput274 output274/A vssd1 vssd1 vccd1 vccd1 y_i_0[7] sky130_fd_sc_hd__buf_2
XFILLER_87_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput285 output285/A vssd1 vssd1 vccd1 vccd1 y_i_1[1] sky130_fd_sc_hd__buf_2
XANTENNA__08160__B _11491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput296 _10934_/X vssd1 vssd1 vccd1 vccd1 y_i_2[11] sky130_fd_sc_hd__buf_2
XFILLER_134_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08940__A2 _15447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _15709_/Q vssd1 vssd1 vccd1 vccd1 _11248_/A sky130_fd_sc_hd__inv_2
XFILLER_210_1123 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09707_ _09699_/Y _09703_/B _09701_/B vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__o21ai_1
X_07899_ _07899_/A vssd1 vssd1 vccd1 vccd1 _15318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09638_ _09636_/A _09636_/B _09637_/X vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07900__A0 _15317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09569_ _15435_/Q _15419_/Q vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14618__A _14620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__S _11928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _12228_/A _11600_/B _11600_/C vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__and3_1
XFILLER_90_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _14940_/Q _12580_/B vssd1 vssd1 vccd1 vccd1 _12580_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11531_ _11531_/A vssd1 vssd1 vccd1 vccd1 _11531_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14250_/Y sky130_fd_sc_hd__inv_2
X_11462_ _11462_/A _11462_/B vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__or2_2
XFILLER_17_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13201_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__or2_1
XANTENNA__11977__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10413_ _10412_/B _10412_/C _10412_/A vssd1 vssd1 vccd1 vccd1 _10417_/B sky130_fd_sc_hd__o21ai_1
X_14181_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14181_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11393_ _15070_/Q _15235_/Q _10191_/Y _09688_/Y vssd1 vssd1 vccd1 vccd1 _11394_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14353__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _13290_/A _13700_/A _13063_/A vssd1 vssd1 vccd1 vccd1 _13133_/B sky130_fd_sc_hd__a21o_1
XFILLER_174_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input62_A x_i_3[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ _10341_/A _10469_/A _10341_/B _10343_/X vssd1 vssd1 vccd1 vccd1 _10347_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08351__A _14938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1048 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _13063_/A _13063_/B vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__nor2_4
X_10275_ _10274_/A _10274_/B _11421_/A vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__a21o_1
XFILLER_79_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _12014_/A _12014_/B vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__xnor2_2
XFILLER_78_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1051 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13416__B _15052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13965_ _13977_/A vssd1 vssd1 vccd1 vccd1 _13965_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output316_A _15674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _15705_/CLK _15704_/D _14779_/Y vssd1 vssd1 vccd1 vccd1 _15704_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_1114 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12916_ _13677_/C _12916_/B vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__xnor2_4
XFILLER_111_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13896_ _08801_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _13897_/C sky130_fd_sc_hd__and2b_1
XFILLER_206_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15635_ _15768_/CLK _15635_/D _14707_/Y vssd1 vssd1 vccd1 vccd1 _15635_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12847_ _15761_/Q vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__inv_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14528__A _14538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _15571_/CLK _15566_/D _14633_/Y vssd1 vssd1 vccd1 vccd1 _15566_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_203_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12771_/A _12776_/X _12771_/B _12777_/X vssd1 vssd1 vccd1 vccd1 _12841_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_148_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10775__B _15786_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14517_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14517_/Y sky130_fd_sc_hd__inv_2
X_11729_ _11651_/A _11651_/B _11718_/X _11728_/Y _11719_/X vssd1 vssd1 vccd1 vccd1
+ _11783_/B sky130_fd_sc_hd__a311oi_4
XFILLER_159_276 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15497_ _15572_/CLK _15497_/D _14560_/Y vssd1 vssd1 vccd1 vccd1 _15497_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ _14460_/A vssd1 vssd1 vccd1 vccd1 _14448_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_repeater800_A repeater801/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14379_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14379_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14263__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1001 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ _15463_/Q _15447_/Q _08939_/B vssd1 vssd1 vccd1 vccd1 _08940_/X sky130_fd_sc_hd__o21a_1
XFILLER_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_891 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ _08947_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _15206_/D sky130_fd_sc_hd__xor2_1
XFILLER_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater700 _07795_/S vssd1 vssd1 vccd1 vccd1 _07803_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07822_ _15356_/Q _07822_/A1 _07856_/S vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__mux2_1
Xrepeater711 _07434_/A vssd1 vssd1 vccd1 vccd1 _07900_/S sky130_fd_sc_hd__buf_6
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12511__A _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__B _15425_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater722 _15693_/Q vssd1 vssd1 vccd1 vccd1 output387/A sky130_fd_sc_hd__clkbuf_2
Xrepeater733 _15675_/Q vssd1 vssd1 vccd1 vccd1 repeater733/X sky130_fd_sc_hd__buf_4
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater744 _15656_/Q vssd1 vssd1 vccd1 vccd1 output281/A sky130_fd_sc_hd__clkbuf_2
Xrepeater755 repeater756/X vssd1 vssd1 vccd1 vccd1 output287/A sky130_fd_sc_hd__buf_6
XANTENNA__09092__A _15499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _15390_/Q _07753_/A1 _07765_/S vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater766 _15633_/Q vssd1 vssd1 vccd1 vccd1 output529/A sky130_fd_sc_hd__clkbuf_2
Xrepeater777 _15620_/Q vssd1 vssd1 vccd1 vccd1 repeater777/X sky130_fd_sc_hd__buf_2
XFILLER_42_1195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater788 _15604_/Q vssd1 vssd1 vccd1 vccd1 repeater788/X sky130_fd_sc_hd__buf_2
Xrepeater799 _15592_/Q vssd1 vssd1 vccd1 vccd1 output419/A sky130_fd_sc_hd__clkbuf_2
X_07684_ _07684_/A vssd1 vssd1 vccd1 vccd1 _15424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_396 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ _09421_/Y _09423_/B vssd1 vssd1 vccd1 vccd1 _09504_/A sky130_fd_sc_hd__nand2b_1
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14438__A _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _09354_/A _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__and3_1
XFILLER_12_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08305_ _08305_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08310_/A sky130_fd_sc_hd__nor2_1
X_09285_ _15400_/Q _15384_/Q vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11993__A1 _12144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08236_ _08292_/B _08236_/B vssd1 vssd1 vccd1 vccd1 _08237_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11797__A _11797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ _15012_/Q vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__buf_6
XANTENNA__07994__B _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14173__A _14176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08098_ _11876_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10060_ _10060_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12170__A1 _12238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10962_ _10962_/A _11143_/A vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_141_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input214_A x_r_5[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ _13849_/B _13849_/C _14981_/Q vssd1 vssd1 vccd1 vccd1 _13752_/A sky130_fd_sc_hd__a21boi_1
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12701_ _12699_/Y _13528_/B _12700_/X vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__o21ai_1
XFILLER_204_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _10891_/Y _10893_/B vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__and2b_1
X_13681_ _13681_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13682_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14348__A _14359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15420_ _15808_/CLK _15420_/D _14479_/Y vssd1 vssd1 vccd1 vccd1 _15420_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12632_ _13203_/A _12945_/A vssd1 vssd1 vccd1 vccd1 _12632_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_34_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12563_ _12563_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _15622_/D sky130_fd_sc_hd__xnor2_1
X_15351_ _15754_/CLK _15351_/D _14406_/Y vssd1 vssd1 vccd1 vccd1 _15351_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1014 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1134 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1088 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ _11898_/A _11797_/A _11587_/B vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__and3_1
XFILLER_12_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14302_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14302_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12494_ _14951_/Q _12504_/B vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__or2_1
X_15282_ _15399_/CLK _15282_/D _14333_/Y vssd1 vssd1 vccd1 vccd1 _15282_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_779 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ _11876_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__nand2_1
X_14233_ _14238_/A vssd1 vssd1 vccd1 vccd1 _14233_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14083__A _14098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07396__S _07432_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _14178_/A vssd1 vssd1 vccd1 vccd1 _14164_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11376_ _11375_/B _11375_/C _11375_/A vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__o21a_1
XFILLER_152_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_963 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _15127_/Q _15160_/Q vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__nor2_1
X_13115_ _13165_/A _13165_/B vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__xnor2_1
XFILLER_180_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14095_ _14098_/A vssd1 vssd1 vccd1 vccd1 _14095_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14811__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _13046_/B vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__or2_1
XFILLER_140_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _15245_/Q _15080_/Q vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__or2b_1
XANTENNA_output433_A output433/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _15070_/Q _15235_/Q vssd1 vssd1 vccd1 vccd1 _10190_/B sky130_fd_sc_hd__or2b_1
XFILLER_67_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater583_A _11197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ _15498_/CLK _14997_/D _14031_/Y vssd1 vssd1 vccd1 vccd1 _14997_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13948_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13948_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13879_ _15335_/Q _15319_/Q _13878_/X vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__a21o_1
XFILLER_61_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14258__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15618_ _15784_/CLK _15618_/D _14689_/Y vssd1 vssd1 vccd1 vccd1 _15618_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_210_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_859 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15549_ _15569_/CLK _15549_/D _14615_/Y vssd1 vssd1 vccd1 vccd1 _15549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09070_ _15493_/Q _15477_/Q _09219_/C vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08021_ _12308_/S _11438_/B vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__xnor2_1
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15239__D _15239_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15817__A _15817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09972_ _15186_/Q _15219_/Q _09869_/Y _10380_/A vssd1 vssd1 vccd1 vccd1 _09973_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14721__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ _08923_/A _08925_/B vssd1 vssd1 vccd1 vccd1 _15214_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_1235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13337__A _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ _15463_/Q _15447_/Q vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__xnor2_1
XFILLER_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _07805_/A vssd1 vssd1 vccd1 vccd1 _07856_/S sky130_fd_sc_hd__buf_12
Xrepeater541 _11296_/X vssd1 vssd1 vccd1 vccd1 output469/A sky130_fd_sc_hd__clkbuf_2
Xrepeater552 _10947_/X vssd1 vssd1 vccd1 vccd1 _10948_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _08783_/Y _08785_/B vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__nand2b_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater563 _11134_/X vssd1 vssd1 vccd1 vccd1 output366/A sky130_fd_sc_hd__buf_4
XFILLER_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater574 _11377_/Y vssd1 vssd1 vccd1 vccd1 output432/A sky130_fd_sc_hd__buf_4
XFILLER_211_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07736_ _15398_/Q input218/X _07750_/S vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__mux2_1
Xrepeater585 _11071_/X vssd1 vssd1 vccd1 vccd1 output262/A sky130_fd_sc_hd__clkbuf_2
Xrepeater596 _11183_/Y vssd1 vssd1 vccd1 vccd1 output511/A sky130_fd_sc_hd__clkbuf_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07667_ _15432_/Q input252/X _07697_/S vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14168__A _14178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1039 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ _15509_/Q vssd1 vssd1 vccd1 vccd1 _09411_/B sky130_fd_sc_hd__inv_2
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08166__A _11906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07598_ _15466_/Q input78/X _07640_/S vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09337_ _15410_/Q _15394_/Q vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09268_ _09268_/A _09268_/B vssd1 vssd1 vccd1 vccd1 _15248_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08219_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__xnor2_2
XFILLER_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09199_ _15573_/Q _15553_/Q vssd1 vssd1 vccd1 vccd1 _09667_/B sky130_fd_sc_hd__xor2_2
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11230_/A _11230_/B _11382_/A vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__and3_1
XFILLER_88_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07398__A1 _07398_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11161_ _11357_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__xor2_1
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input164_A x_r_2[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14631__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10112_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__nand2_2
XANTENNA__09139__A2 _15491_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11348_/A sky130_fd_sc_hd__nor2_2
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ _10043_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14920_ _15532_/CLK _14920_/D _13950_/Y vssd1 vssd1 vccd1 vccd1 _14920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_79 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_707 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12151__A _12466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14851_ _14853_/A vssd1 vssd1 vccd1 vccd1 _14851_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input25_A x_i_1[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13791_/A _13791_/B _13801_/X vssd1 vssd1 vccd1 vccd1 _13806_/A sky130_fd_sc_hd__a21o_1
XFILLER_5_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__buf_6
XFILLER_112_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _11912_/A _11994_/B _11994_/C vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__and3b_1
XFILLER_21_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10457__A1 _15125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ _13721_/A _13832_/B _13838_/B _13732_/Y _13728_/A vssd1 vssd1 vccd1 vccd1
+ _13743_/A sky130_fd_sc_hd__o311a_1
XFILLER_189_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10945_ _10945_/A _10945_/B _11134_/A vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__and3_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14078__A _14078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15612__D _15612_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _13815_/A _13664_/B vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__xnor2_4
X_10876_ _11109_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10881_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ _15406_/CLK _15403_/D _14462_/Y vssd1 vssd1 vccd1 vccd1 _15403_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _14952_/Q vssd1 vssd1 vccd1 vccd1 _12615_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13595_ _15367_/Q _15351_/Q _13594_/B vssd1 vssd1 vccd1 vccd1 _13595_/X sky130_fd_sc_hd__o21a_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14806__A _14821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15428_/CLK _15334_/D _14388_/Y vssd1 vssd1 vccd1 vccd1 _15334_/Q sky130_fd_sc_hd__dfrtp_1
X_12546_ _12543_/A _12544_/A _12543_/B _12545_/X vssd1 vssd1 vccd1 vccd1 _12548_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA_output383_A output383/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15265_ _15539_/CLK _15265_/D _14315_/Y vssd1 vssd1 vccd1 vccd1 _15265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _12601_/A _12604_/A vssd1 vssd1 vccd1 vccd1 _12478_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14216_ _14218_/A vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__inv_2
X_11428_ _15084_/Q _15249_/Q vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_1221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15196_ _15472_/CLK _15196_/D _14243_/Y vssd1 vssd1 vccd1 vccd1 _15196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11359_/Y sky130_fd_sc_hd__xnor2_2
X_14147_ _14158_/A vssd1 vssd1 vccd1 vccd1 _14147_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07854__S _07856_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14078_ _14078_/A vssd1 vssd1 vccd1 vccd1 _14078_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater798_A _15593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1015 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ _13162_/B _13102_/B vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13882__A1 _15336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_564 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1025 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07561__A1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08570_ _08570_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07521_ _07521_/A vssd1 vssd1 vccd1 vccd1 _15504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07452_ _07452_/A vssd1 vssd1 vccd1 vccd1 _15538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13323__C _13381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _07383_/A vssd1 vssd1 vccd1 vccd1 _15576_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14716__A _14721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ _15504_/Q _15488_/Q vssd1 vssd1 vccd1 vccd1 _09122_/X sky130_fd_sc_hd__and2_1
XFILLER_175_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ _09052_/A _09052_/B _13625_/A vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__a21oi_1
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ _08004_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__xor2_1
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_719 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14451__A _14460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _09953_/X _09958_/B vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08906_ _08906_/A _08914_/A vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__nand2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _15189_/Q _15222_/Q vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__nand2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ _08836_/A _08836_/B _13911_/A vssd1 vssd1 vccd1 vccd1 _08838_/B sky130_fd_sc_hd__o21a_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08768_ _08768_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _15071_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_439 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _07719_/A vssd1 vssd1 vccd1 vccd1 _15407_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08699_ _08699_/A _12692_/B vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__xnor2_4
XFILLER_54_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08608__B _12803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10730_ _15712_/Q _15778_/Q vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ _15274_/Q _15175_/Q vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14626__A _14640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12400_ _12400_/A vssd1 vssd1 vccd1 vccd1 _15648_/D sky130_fd_sc_hd__clkbuf_1
X_13380_ _13380_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _13384_/A sky130_fd_sc_hd__xnor2_1
XFILLER_210_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10592_ _10592_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _14989_/D sky130_fd_sc_hd__xnor2_1
XFILLER_107_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _12331_/A vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__inv_2
XFILLER_103_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12262_ _12262_/A _12491_/A vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__or2_1
X_15050_ _15693_/CLK _15050_/D _14088_/Y vssd1 vssd1 vccd1 vccd1 _15050_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14001_ _14003_/A vssd1 vssd1 vccd1 vccd1 _14001_/Y sky130_fd_sc_hd__inv_2
X_11213_ _15753_/Q _15031_/Q vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__or2b_1
X_12193_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12194_/B sky130_fd_sc_hd__and2_1
XANTENNA__14361__A _14369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11144_ _15021_/Q _15743_/Q vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__or2b_1
XANTENNA__09780__A2 _15416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_989 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07791__A1 input239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11075_ _14999_/Q _14933_/Q vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__and2b_1
XFILLER_122_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput130 x_i_7[9] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput141 x_r_0[4] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__clkbuf_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10678__A1 _15276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14903_ _15732_/CLK _14903_/D _13932_/Y vssd1 vssd1 vccd1 vccd1 _14903_/Q sky130_fd_sc_hd__dfrtp_1
X_10026_ _15205_/Q _15106_/Q vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__nor2_1
Xinput152 x_r_1[14] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_4
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput163 x_r_2[0] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__clkbuf_1
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput174 x_r_2[5] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07543__A1 _07543_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput185 x_r_3[15] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_4
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 x_r_4[10] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__buf_4
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _14836_/A vssd1 vssd1 vccd1 vccd1 _14834_/Y sky130_fd_sc_hd__inv_2
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _14774_/A vssd1 vssd1 vccd1 vccd1 _14765_/Y sky130_fd_sc_hd__inv_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11977_ _11977_/A _11977_/B vssd1 vssd1 vccd1 vccd1 _11978_/B sky130_fd_sc_hd__or2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13716_ _13725_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__nand2_1
X_10928_ _14965_/Q _14899_/Q vssd1 vssd1 vccd1 vccd1 _10930_/A sky130_fd_sc_hd__or2b_1
X_14696_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14696_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13647_ _13669_/A _13646_/B _13646_/C vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__a21o_1
X_10859_ _10867_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__nand2_1
XANTENNA_repeater546_A _12575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_829 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14536__A _14540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11879__B _12231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08534__A _08728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ _13574_/A _13571_/A _13577_/X vssd1 vssd1 vccd1 vccd1 _13579_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10783__B _15787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ _15722_/CLK _15317_/D _14370_/Y vssd1 vssd1 vccd1 vccd1 _15317_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_8_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ _12529_/A _12529_/B vssd1 vssd1 vccd1 vccd1 _15612_/D sky130_fd_sc_hd__xnor2_1
XFILLER_157_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater713_A _15707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_885 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15248_ _15347_/CLK _15248_/D _14297_/Y vssd1 vssd1 vccd1 vccd1 _15248_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_207_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15179_ _15180_/CLK _15179_/D _14224_/Y vssd1 vssd1 vccd1 vccd1 _15179_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14271__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1122 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1027 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1035 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09740_ _15064_/Q _15097_/Q vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

